magic
tech sky130A
timestamp 1697129952
<< nwell >>
rect -115 695 1675 2060
<< nmos >>
rect 5 -20 55 580
rect 105 -20 155 580
rect 205 -20 255 580
rect 305 -20 355 580
rect 405 -20 455 580
rect 505 -20 555 580
rect 605 -20 655 580
rect 705 -20 755 580
rect 805 -20 855 580
rect 905 -20 955 580
rect 1005 -20 1055 580
rect 1105 -20 1155 580
rect 1205 -20 1255 580
rect 1305 -20 1355 580
rect 1405 -20 1455 580
rect 1505 -20 1555 580
rect 5 -745 55 -145
rect 105 -745 155 -145
rect 205 -745 255 -145
rect 305 -745 355 -145
rect 405 -745 455 -145
rect 505 -745 555 -145
rect 605 -745 655 -145
rect 705 -745 755 -145
rect 805 -745 855 -145
rect 905 -745 955 -145
rect 1005 -745 1055 -145
rect 1105 -745 1155 -145
rect 1205 -745 1255 -145
rect 1305 -745 1355 -145
rect 1405 -745 1455 -145
rect 1505 -745 1555 -145
<< pmos >>
rect 5 1440 55 2040
rect 105 1440 155 2040
rect 205 1440 255 2040
rect 305 1440 355 2040
rect 405 1440 455 2040
rect 505 1440 555 2040
rect 605 1440 655 2040
rect 705 1440 755 2040
rect 805 1440 855 2040
rect 905 1440 955 2040
rect 1005 1440 1055 2040
rect 1105 1440 1155 2040
rect 1205 1440 1255 2040
rect 1305 1440 1355 2040
rect 1405 1440 1455 2040
rect 1505 1440 1555 2040
rect 5 715 55 1315
rect 105 715 155 1315
rect 205 715 255 1315
rect 305 715 355 1315
rect 405 715 455 1315
rect 505 715 555 1315
rect 605 715 655 1315
rect 705 715 755 1315
rect 805 715 855 1315
rect 905 715 955 1315
rect 1005 715 1055 1315
rect 1105 715 1155 1315
rect 1205 715 1255 1315
rect 1305 715 1355 1315
rect 1405 715 1455 1315
rect 1505 715 1555 1315
<< ndiff >>
rect -45 565 5 580
rect -45 -5 -30 565
rect -10 -5 5 565
rect -45 -20 5 -5
rect 55 565 105 580
rect 55 -5 70 565
rect 90 -5 105 565
rect 55 -20 105 -5
rect 155 565 205 580
rect 155 -5 170 565
rect 190 -5 205 565
rect 155 -20 205 -5
rect 255 565 305 580
rect 255 -5 270 565
rect 290 -5 305 565
rect 255 -20 305 -5
rect 355 565 405 580
rect 355 -5 370 565
rect 390 -5 405 565
rect 355 -20 405 -5
rect 455 565 505 580
rect 455 -5 470 565
rect 490 -5 505 565
rect 455 -20 505 -5
rect 555 565 605 580
rect 555 -5 570 565
rect 590 -5 605 565
rect 555 -20 605 -5
rect 655 565 705 580
rect 655 -5 670 565
rect 690 -5 705 565
rect 655 -20 705 -5
rect 755 565 805 580
rect 755 -5 770 565
rect 790 -5 805 565
rect 755 -20 805 -5
rect 855 565 905 580
rect 855 -5 870 565
rect 890 -5 905 565
rect 855 -20 905 -5
rect 955 565 1005 580
rect 955 -5 970 565
rect 990 -5 1005 565
rect 955 -20 1005 -5
rect 1055 565 1105 580
rect 1055 -5 1070 565
rect 1090 -5 1105 565
rect 1055 -20 1105 -5
rect 1155 565 1205 580
rect 1155 -5 1170 565
rect 1190 -5 1205 565
rect 1155 -20 1205 -5
rect 1255 565 1305 580
rect 1255 -5 1270 565
rect 1290 -5 1305 565
rect 1255 -20 1305 -5
rect 1355 565 1405 580
rect 1355 -5 1370 565
rect 1390 -5 1405 565
rect 1355 -20 1405 -5
rect 1455 565 1505 580
rect 1455 -5 1470 565
rect 1490 -5 1505 565
rect 1455 -20 1505 -5
rect 1555 565 1605 580
rect 1555 -5 1570 565
rect 1590 -5 1605 565
rect 1555 -20 1605 -5
rect -45 -160 5 -145
rect -45 -730 -30 -160
rect -10 -730 5 -160
rect -45 -745 5 -730
rect 55 -160 105 -145
rect 55 -730 70 -160
rect 90 -730 105 -160
rect 55 -745 105 -730
rect 155 -160 205 -145
rect 155 -730 170 -160
rect 190 -730 205 -160
rect 155 -745 205 -730
rect 255 -745 305 -145
rect 355 -745 405 -145
rect 455 -745 505 -145
rect 555 -745 605 -145
rect 655 -745 705 -145
rect 755 -160 805 -145
rect 755 -730 770 -160
rect 790 -730 805 -160
rect 755 -745 805 -730
rect 855 -745 905 -145
rect 955 -745 1005 -145
rect 1055 -745 1105 -145
rect 1155 -745 1205 -145
rect 1255 -745 1305 -145
rect 1355 -160 1405 -145
rect 1355 -730 1370 -160
rect 1390 -730 1405 -160
rect 1355 -745 1405 -730
rect 1455 -160 1505 -145
rect 1455 -730 1470 -160
rect 1490 -730 1505 -160
rect 1455 -745 1505 -730
rect 1555 -160 1605 -145
rect 1555 -730 1570 -160
rect 1590 -730 1605 -160
rect 1555 -745 1605 -730
<< pdiff >>
rect -45 2025 5 2040
rect -45 1455 -30 2025
rect -10 1455 5 2025
rect -45 1440 5 1455
rect 55 2025 105 2040
rect 55 1455 70 2025
rect 90 1455 105 2025
rect 55 1440 105 1455
rect 155 2025 205 2040
rect 155 1455 170 2025
rect 190 1455 205 2025
rect 155 1440 205 1455
rect 255 1440 305 2040
rect 355 1440 405 2040
rect 455 1440 505 2040
rect 555 1440 605 2040
rect 655 1440 705 2040
rect 755 2025 805 2040
rect 755 1455 770 2025
rect 790 1455 805 2025
rect 755 1440 805 1455
rect 855 1440 905 2040
rect 955 1440 1005 2040
rect 1055 1440 1105 2040
rect 1155 1440 1205 2040
rect 1255 1440 1305 2040
rect 1355 2025 1405 2040
rect 1355 1455 1370 2025
rect 1390 1455 1405 2025
rect 1355 1440 1405 1455
rect 1455 2025 1505 2040
rect 1455 1455 1470 2025
rect 1490 1455 1505 2025
rect 1455 1440 1505 1455
rect 1555 2025 1605 2040
rect 1555 1455 1570 2025
rect 1590 1455 1605 2025
rect 1555 1440 1605 1455
rect -45 1300 5 1315
rect -45 730 -30 1300
rect -10 730 5 1300
rect -45 715 5 730
rect 55 1300 105 1315
rect 55 730 70 1300
rect 90 730 105 1300
rect 55 715 105 730
rect 155 1300 205 1315
rect 155 730 170 1300
rect 190 730 205 1300
rect 155 715 205 730
rect 255 1300 305 1315
rect 255 730 270 1300
rect 290 730 305 1300
rect 255 715 305 730
rect 355 1300 405 1315
rect 355 730 370 1300
rect 390 730 405 1300
rect 355 715 405 730
rect 455 1300 505 1315
rect 455 730 470 1300
rect 490 730 505 1300
rect 455 715 505 730
rect 555 1300 605 1315
rect 555 730 570 1300
rect 590 730 605 1300
rect 555 715 605 730
rect 655 1300 705 1315
rect 655 730 670 1300
rect 690 730 705 1300
rect 655 715 705 730
rect 755 1300 805 1315
rect 755 730 770 1300
rect 790 730 805 1300
rect 755 715 805 730
rect 855 1300 905 1315
rect 855 730 870 1300
rect 890 730 905 1300
rect 855 715 905 730
rect 955 1300 1005 1315
rect 955 730 970 1300
rect 990 730 1005 1300
rect 955 715 1005 730
rect 1055 1300 1105 1315
rect 1055 730 1070 1300
rect 1090 730 1105 1300
rect 1055 715 1105 730
rect 1155 1300 1205 1315
rect 1155 730 1170 1300
rect 1190 730 1205 1300
rect 1155 715 1205 730
rect 1255 1300 1305 1315
rect 1255 730 1270 1300
rect 1290 730 1305 1300
rect 1255 715 1305 730
rect 1355 1300 1405 1315
rect 1355 730 1370 1300
rect 1390 730 1405 1300
rect 1355 715 1405 730
rect 1455 1300 1505 1315
rect 1455 730 1470 1300
rect 1490 730 1505 1300
rect 1455 715 1505 730
rect 1555 1300 1605 1315
rect 1555 730 1570 1300
rect 1590 730 1605 1300
rect 1555 715 1605 730
<< ndiffc >>
rect -30 -5 -10 565
rect 70 -5 90 565
rect 170 -5 190 565
rect 270 -5 290 565
rect 370 -5 390 565
rect 470 -5 490 565
rect 570 -5 590 565
rect 670 -5 690 565
rect 770 -5 790 565
rect 870 -5 890 565
rect 970 -5 990 565
rect 1070 -5 1090 565
rect 1170 -5 1190 565
rect 1270 -5 1290 565
rect 1370 -5 1390 565
rect 1470 -5 1490 565
rect 1570 -5 1590 565
rect -30 -730 -10 -160
rect 70 -730 90 -160
rect 170 -730 190 -160
rect 770 -730 790 -160
rect 1370 -730 1390 -160
rect 1470 -730 1490 -160
rect 1570 -730 1590 -160
<< pdiffc >>
rect -30 1455 -10 2025
rect 70 1455 90 2025
rect 170 1455 190 2025
rect 770 1455 790 2025
rect 1370 1455 1390 2025
rect 1470 1455 1490 2025
rect 1570 1455 1590 2025
rect -30 730 -10 1300
rect 70 730 90 1300
rect 170 730 190 1300
rect 270 730 290 1300
rect 370 730 390 1300
rect 470 730 490 1300
rect 570 730 590 1300
rect 670 730 690 1300
rect 770 730 790 1300
rect 870 730 890 1300
rect 970 730 990 1300
rect 1070 730 1090 1300
rect 1170 730 1190 1300
rect 1270 730 1290 1300
rect 1370 730 1390 1300
rect 1470 730 1490 1300
rect 1570 730 1590 1300
<< psubdiff >>
rect -95 565 -45 580
rect -95 -5 -80 565
rect -60 -5 -45 565
rect -95 -20 -45 -5
rect 1605 565 1655 580
rect 1605 -5 1620 565
rect 1640 -5 1655 565
rect 1605 -20 1655 -5
rect -95 -160 -45 -145
rect -95 -730 -80 -160
rect -60 -730 -45 -160
rect -95 -745 -45 -730
rect 1605 -160 1655 -145
rect 1605 -730 1620 -160
rect 1640 -730 1655 -160
rect 1605 -745 1655 -730
<< nsubdiff >>
rect -95 2025 -45 2040
rect -95 1455 -80 2025
rect -60 1455 -45 2025
rect -95 1440 -45 1455
rect 1605 2025 1655 2040
rect 1605 1455 1620 2025
rect 1640 1455 1655 2025
rect 1605 1440 1655 1455
rect -95 1300 -45 1315
rect -95 730 -80 1300
rect -60 730 -45 1300
rect -95 715 -45 730
rect 1605 1300 1655 1315
rect 1605 730 1620 1300
rect 1640 730 1655 1300
rect 1605 715 1655 730
<< psubdiffcont >>
rect -80 -5 -60 565
rect 1620 -5 1640 565
rect -80 -730 -60 -160
rect 1620 -730 1640 -160
<< nsubdiffcont >>
rect -80 1455 -60 2025
rect 1620 1455 1640 2025
rect -80 730 -60 1300
rect 1620 730 1640 1300
<< poly >>
rect 1410 2080 1655 2095
rect 1410 2065 1455 2080
rect 5 2040 55 2055
rect 105 2050 1455 2065
rect 105 2040 155 2050
rect 205 2040 255 2050
rect 305 2040 355 2050
rect 405 2040 455 2050
rect 505 2040 555 2050
rect 605 2040 655 2050
rect 705 2040 755 2050
rect 805 2040 855 2050
rect 905 2040 955 2050
rect 1005 2040 1055 2050
rect 1105 2040 1155 2050
rect 1205 2040 1255 2050
rect 1305 2040 1355 2050
rect 1405 2040 1455 2050
rect 1505 2040 1555 2055
rect 5 1425 55 1440
rect 105 1425 155 1440
rect 205 1425 255 1440
rect 305 1425 355 1440
rect 405 1425 455 1440
rect 505 1425 555 1440
rect 605 1425 655 1440
rect -40 1415 55 1425
rect -40 1395 -30 1415
rect -10 1410 55 1415
rect 705 1415 755 1440
rect 805 1415 855 1440
rect 905 1425 955 1440
rect 1005 1425 1055 1440
rect 1105 1425 1155 1440
rect 1205 1425 1255 1440
rect 1305 1425 1355 1440
rect 1405 1425 1455 1440
rect 1505 1425 1555 1440
rect -10 1395 0 1410
rect -40 1385 0 1395
rect 705 1405 855 1415
rect 1505 1415 1655 1425
rect 1505 1410 1625 1415
rect 705 1385 770 1405
rect 790 1385 855 1405
rect 1615 1395 1625 1410
rect 1645 1395 1655 1415
rect 1615 1385 1655 1395
rect 705 1375 855 1385
rect 5 1315 55 1330
rect 105 1315 155 1330
rect 205 1315 255 1330
rect 305 1315 355 1330
rect 405 1315 455 1330
rect 505 1315 555 1330
rect 605 1315 655 1330
rect 705 1315 755 1375
rect 805 1315 855 1375
rect 1405 1355 1590 1370
rect 905 1315 955 1330
rect 1005 1315 1055 1330
rect 1105 1315 1155 1330
rect 1205 1315 1255 1330
rect 1305 1315 1355 1330
rect 1405 1315 1455 1355
rect 1575 1340 1655 1355
rect 1505 1315 1555 1330
rect 5 700 55 715
rect -40 690 55 700
rect -40 670 -30 690
rect -10 685 55 690
rect 105 690 155 715
rect -10 670 0 685
rect -40 660 0 670
rect 105 670 120 690
rect 140 670 155 690
rect 105 660 155 670
rect 205 690 255 715
rect 205 670 220 690
rect 240 670 255 690
rect 205 660 255 670
rect 305 690 355 715
rect 305 670 320 690
rect 340 670 355 690
rect 305 660 355 670
rect 405 690 455 715
rect 405 670 420 690
rect 440 670 455 690
rect 405 660 455 670
rect 505 690 555 715
rect 505 670 520 690
rect 540 670 555 690
rect 505 660 555 670
rect 605 690 655 715
rect 705 700 755 715
rect 805 700 855 715
rect 605 670 620 690
rect 640 670 655 690
rect 605 660 655 670
rect 905 690 955 715
rect 905 670 920 690
rect 940 670 955 690
rect 905 660 955 670
rect 1005 690 1055 715
rect 1005 670 1020 690
rect 1040 670 1055 690
rect 1005 660 1055 670
rect 1105 690 1155 715
rect 1105 670 1120 690
rect 1140 670 1155 690
rect 1105 660 1155 670
rect 1205 690 1255 715
rect 1205 670 1220 690
rect 1240 670 1255 690
rect 1205 660 1255 670
rect 1305 690 1355 715
rect 1305 670 1320 690
rect 1340 670 1355 690
rect 1305 660 1355 670
rect 1405 690 1455 715
rect 1405 670 1420 690
rect 1440 670 1455 690
rect 1505 700 1555 715
rect 1505 690 1600 700
rect 1505 685 1570 690
rect 1405 660 1455 670
rect 1560 670 1570 685
rect 1590 670 1600 690
rect 1560 660 1600 670
rect -40 625 0 635
rect -40 605 -30 625
rect -10 610 0 625
rect 105 625 155 635
rect -10 605 55 610
rect -40 595 55 605
rect 5 580 55 595
rect 105 605 120 625
rect 140 605 155 625
rect 105 580 155 605
rect 205 625 255 635
rect 205 605 220 625
rect 240 605 255 625
rect 205 580 255 605
rect 305 625 355 635
rect 305 605 320 625
rect 340 605 355 625
rect 305 580 355 605
rect 405 625 455 635
rect 405 605 420 625
rect 440 605 455 625
rect 405 580 455 605
rect 505 625 555 635
rect 505 605 520 625
rect 540 605 555 625
rect 505 580 555 605
rect 605 625 655 635
rect 605 605 620 625
rect 640 605 655 625
rect 605 580 655 605
rect 905 625 955 635
rect 905 605 920 625
rect 940 605 955 625
rect 705 580 755 595
rect 805 580 855 595
rect 905 580 955 605
rect 1005 625 1055 635
rect 1005 605 1020 625
rect 1040 605 1055 625
rect 1005 580 1055 605
rect 1105 625 1155 635
rect 1105 605 1120 625
rect 1140 605 1155 625
rect 1105 580 1155 605
rect 1205 625 1255 635
rect 1205 605 1220 625
rect 1240 605 1255 625
rect 1205 580 1255 605
rect 1305 625 1355 635
rect 1305 605 1320 625
rect 1340 605 1355 625
rect 1305 580 1355 605
rect 1405 625 1455 635
rect 1405 605 1420 625
rect 1440 605 1455 625
rect 1560 625 1600 635
rect 1560 610 1570 625
rect 1405 580 1455 605
rect 1505 605 1570 610
rect 1590 605 1600 625
rect 1505 595 1600 605
rect 1505 580 1555 595
rect 5 -35 55 -20
rect 105 -35 155 -20
rect 205 -35 255 -20
rect 305 -35 355 -20
rect 405 -35 455 -20
rect 505 -35 555 -20
rect 605 -35 655 -20
rect -40 -100 0 -90
rect -40 -120 -30 -100
rect -10 -115 0 -100
rect -10 -120 55 -115
rect -40 -130 55 -120
rect 5 -145 55 -130
rect 105 -145 155 -130
rect 205 -145 255 -130
rect 305 -145 355 -130
rect 405 -145 455 -130
rect 505 -145 555 -130
rect 605 -145 655 -130
rect 705 -145 755 -20
rect 805 -145 855 -20
rect 905 -35 955 -20
rect 1005 -35 1055 -20
rect 1105 -35 1155 -20
rect 1205 -35 1255 -20
rect 1305 -35 1355 -20
rect 1405 -60 1455 -20
rect 1505 -35 1555 -20
rect 1580 -60 1655 -45
rect 1405 -75 1595 -60
rect 1615 -100 1655 -90
rect 1615 -115 1625 -100
rect 1505 -120 1625 -115
rect 1645 -120 1655 -100
rect 1505 -130 1655 -120
rect 905 -145 955 -130
rect 1005 -145 1055 -130
rect 1105 -145 1155 -130
rect 1205 -145 1255 -130
rect 1305 -145 1355 -130
rect 1405 -145 1455 -130
rect 1505 -145 1555 -130
rect 5 -760 55 -745
rect 105 -755 155 -745
rect 205 -755 255 -745
rect 305 -755 355 -745
rect 405 -755 455 -745
rect 505 -755 555 -745
rect 605 -755 655 -745
rect 705 -755 755 -745
rect 805 -755 855 -745
rect 905 -755 955 -745
rect 1005 -755 1055 -745
rect 1105 -755 1155 -745
rect 1205 -755 1255 -745
rect 1305 -755 1355 -745
rect 1405 -755 1455 -745
rect 105 -770 1455 -755
rect 1505 -760 1555 -745
rect 1410 -785 1455 -770
rect 1410 -800 1655 -785
<< polycont >>
rect -30 1395 -10 1415
rect 770 1385 790 1405
rect 1625 1395 1645 1415
rect -30 670 -10 690
rect 120 670 140 690
rect 220 670 240 690
rect 320 670 340 690
rect 420 670 440 690
rect 520 670 540 690
rect 620 670 640 690
rect 920 670 940 690
rect 1020 670 1040 690
rect 1120 670 1140 690
rect 1220 670 1240 690
rect 1320 670 1340 690
rect 1420 670 1440 690
rect 1570 670 1590 690
rect -30 605 -10 625
rect 120 605 140 625
rect 220 605 240 625
rect 320 605 340 625
rect 420 605 440 625
rect 520 605 540 625
rect 620 605 640 625
rect 920 605 940 625
rect 1020 605 1040 625
rect 1120 605 1140 625
rect 1220 605 1240 625
rect 1320 605 1340 625
rect 1420 605 1440 625
rect 1570 605 1590 625
rect -30 -120 -10 -100
rect 1625 -120 1645 -100
<< locali >>
rect 60 2055 1500 2095
rect -90 2025 0 2035
rect -90 1455 -80 2025
rect -60 1455 -30 2025
rect -10 1455 0 2025
rect -90 1445 0 1455
rect -40 1415 0 1445
rect -40 1395 -30 1415
rect -10 1395 0 1415
rect -40 1385 0 1395
rect 60 2025 100 2055
rect 60 1455 70 2025
rect 90 1455 100 2025
rect 60 1375 100 1455
rect 160 2025 200 2035
rect 160 1455 170 2025
rect 190 1455 200 2025
rect 160 1445 200 1455
rect 760 2025 800 2035
rect 760 1455 770 2025
rect 790 1485 800 2025
rect 1360 2025 1400 2035
rect 790 1455 1055 1485
rect 760 1445 1055 1455
rect 1360 1455 1370 2025
rect 1390 1455 1400 2025
rect 1360 1445 1400 1455
rect 1460 2025 1500 2055
rect 1460 1455 1470 2025
rect 1490 1455 1500 2025
rect 760 1405 800 1415
rect 760 1385 770 1405
rect 790 1385 800 1405
rect 760 1375 800 1385
rect 1005 1405 1055 1445
rect 1005 1385 1015 1405
rect 1045 1385 1055 1405
rect 1005 1375 1055 1385
rect 1460 1375 1500 1455
rect 1560 2025 1650 2035
rect 1560 1455 1570 2025
rect 1590 1455 1620 2025
rect 1640 1455 1650 2025
rect 1560 1445 1650 1455
rect 1615 1425 1650 1445
rect 1615 1415 1655 1425
rect 1615 1395 1625 1415
rect 1645 1395 1655 1415
rect 1615 1385 1655 1395
rect 30 1365 100 1375
rect 30 1345 40 1365
rect 90 1345 100 1365
rect 1460 1365 1530 1375
rect 30 1335 100 1345
rect 160 1335 1400 1355
rect 1460 1345 1470 1365
rect 1520 1345 1530 1365
rect 1460 1335 1530 1345
rect -90 1300 0 1310
rect -90 730 -80 1300
rect -60 730 -30 1300
rect -10 730 0 1300
rect -90 720 0 730
rect -40 690 0 720
rect -40 670 -30 690
rect -10 670 0 690
rect -40 660 0 670
rect 60 1300 100 1310
rect 60 730 70 1300
rect 90 730 100 1300
rect 60 700 100 730
rect 160 1300 200 1335
rect 160 730 170 1300
rect 190 730 200 1300
rect 160 720 200 730
rect 260 1300 300 1310
rect 260 730 270 1300
rect 290 730 300 1300
rect 260 700 300 730
rect 360 1300 400 1335
rect 360 730 370 1300
rect 390 730 400 1300
rect 360 720 400 730
rect 460 1300 500 1310
rect 460 730 470 1300
rect 490 730 500 1300
rect 460 700 500 730
rect 560 1300 600 1335
rect 560 730 570 1300
rect 590 730 600 1300
rect 560 720 600 730
rect 660 1300 700 1310
rect 660 730 670 1300
rect 690 730 700 1300
rect 660 720 700 730
rect 760 1300 800 1310
rect 760 730 770 1300
rect 790 730 800 1300
rect 760 720 800 730
rect 860 1300 900 1310
rect 860 730 870 1300
rect 890 730 900 1300
rect 860 720 900 730
rect 960 1300 1000 1335
rect 960 730 970 1300
rect 990 730 1000 1300
rect 960 720 1000 730
rect 1060 1300 1100 1310
rect 1060 730 1070 1300
rect 1090 730 1100 1300
rect 1060 700 1100 730
rect 1160 1300 1200 1335
rect 1160 730 1170 1300
rect 1190 730 1200 1300
rect 1160 720 1200 730
rect 1260 1300 1300 1310
rect 1260 730 1270 1300
rect 1290 730 1300 1300
rect 1260 700 1300 730
rect 1360 1300 1400 1335
rect 1360 730 1370 1300
rect 1390 730 1400 1300
rect 1360 720 1400 730
rect 1460 1300 1500 1310
rect 1460 730 1470 1300
rect 1490 730 1500 1300
rect 1460 700 1500 730
rect 60 690 155 700
rect 60 670 120 690
rect 140 670 155 690
rect 60 660 155 670
rect 205 690 1355 700
rect 205 670 220 690
rect 240 670 320 690
rect 340 670 420 690
rect 440 670 520 690
rect 540 670 620 690
rect 640 670 920 690
rect 940 670 1020 690
rect 1040 670 1120 690
rect 1140 670 1220 690
rect 1240 670 1320 690
rect 1340 670 1355 690
rect 205 660 1355 670
rect 1405 690 1500 700
rect 1405 670 1420 690
rect 1440 670 1500 690
rect 1405 660 1500 670
rect 1560 1300 1650 1310
rect 1560 730 1570 1300
rect 1590 730 1620 1300
rect 1640 730 1650 1300
rect 1560 720 1650 730
rect 1560 690 1600 720
rect 1560 670 1570 690
rect 1590 670 1600 690
rect 1560 660 1600 670
rect -40 625 0 635
rect -40 605 -30 625
rect -10 605 0 625
rect -40 575 0 605
rect -90 565 0 575
rect -90 -5 -80 565
rect -60 -5 -30 565
rect -10 -5 0 565
rect -90 -15 0 -5
rect 60 625 155 635
rect 60 605 120 625
rect 140 605 155 625
rect 60 595 155 605
rect 205 625 1355 635
rect 205 605 220 625
rect 240 605 320 625
rect 340 605 420 625
rect 440 605 520 625
rect 540 605 620 625
rect 640 605 920 625
rect 940 605 1020 625
rect 1040 605 1120 625
rect 1140 605 1220 625
rect 1240 605 1320 625
rect 1340 605 1355 625
rect 205 595 1355 605
rect 1405 625 1500 635
rect 1405 605 1420 625
rect 1440 605 1500 625
rect 1405 595 1500 605
rect 60 565 100 595
rect 60 -5 70 565
rect 90 -5 100 565
rect 60 -15 100 -5
rect 160 565 200 575
rect 160 -5 170 565
rect 190 -5 200 565
rect 160 -40 200 -5
rect 260 565 300 595
rect 260 -5 270 565
rect 290 -5 300 565
rect 260 -15 300 -5
rect 360 565 400 575
rect 360 -5 370 565
rect 390 -5 400 565
rect 360 -40 400 -5
rect 460 565 500 595
rect 460 -5 470 565
rect 490 -5 500 565
rect 460 -15 500 -5
rect 560 565 600 575
rect 560 -5 570 565
rect 590 -5 600 565
rect 560 -40 600 -5
rect 660 565 700 575
rect 660 -5 670 565
rect 690 -5 700 565
rect 660 -15 700 -5
rect 760 565 800 575
rect 760 -5 770 565
rect 790 -5 800 565
rect 760 -15 800 -5
rect 860 565 900 575
rect 860 -5 870 565
rect 890 -5 900 565
rect 860 -15 900 -5
rect 960 565 1000 575
rect 960 -5 970 565
rect 990 -5 1000 565
rect 960 -40 1000 -5
rect 1060 565 1100 595
rect 1060 -5 1070 565
rect 1090 -5 1100 565
rect 1060 -15 1100 -5
rect 1160 565 1200 575
rect 1160 -5 1170 565
rect 1190 -5 1200 565
rect 1160 -40 1200 -5
rect 1260 565 1300 595
rect 1260 -5 1270 565
rect 1290 -5 1300 565
rect 1260 -15 1300 -5
rect 1360 565 1400 575
rect 1360 -5 1370 565
rect 1390 -5 1400 565
rect 1360 -40 1400 -5
rect 1460 565 1500 595
rect 1460 -5 1470 565
rect 1490 -5 1500 565
rect 1460 -15 1500 -5
rect 1560 625 1600 635
rect 1560 605 1570 625
rect 1590 605 1600 625
rect 1560 575 1600 605
rect 1560 565 1650 575
rect 1560 -5 1570 565
rect 1590 -5 1620 565
rect 1640 -5 1650 565
rect 1560 -15 1650 -5
rect 160 -60 1400 -40
rect 60 -90 255 -80
rect -40 -100 0 -90
rect -40 -120 -30 -100
rect -10 -120 0 -100
rect -40 -150 0 -120
rect -90 -160 0 -150
rect -90 -730 -80 -160
rect -60 -730 -30 -160
rect -10 -730 0 -160
rect -90 -740 0 -730
rect 60 -110 215 -90
rect 245 -110 255 -90
rect 60 -120 255 -110
rect 505 -90 555 -80
rect 505 -110 515 -90
rect 545 -110 555 -90
rect 60 -160 100 -120
rect 505 -150 555 -110
rect 1305 -90 1500 -80
rect 1305 -110 1315 -90
rect 1345 -110 1500 -90
rect 1305 -120 1500 -110
rect 60 -730 70 -160
rect 90 -730 100 -160
rect 60 -760 100 -730
rect 160 -160 200 -150
rect 160 -730 170 -160
rect 190 -730 200 -160
rect 505 -160 800 -150
rect 505 -190 770 -160
rect 160 -740 200 -730
rect 760 -730 770 -190
rect 790 -730 800 -160
rect 760 -740 800 -730
rect 1360 -160 1400 -150
rect 1360 -730 1370 -160
rect 1390 -730 1400 -160
rect 1360 -740 1400 -730
rect 1460 -160 1500 -120
rect 1615 -100 1655 -90
rect 1615 -120 1625 -100
rect 1645 -120 1655 -100
rect 1615 -130 1655 -120
rect 1615 -150 1650 -130
rect 1460 -730 1470 -160
rect 1490 -730 1500 -160
rect 1460 -760 1500 -730
rect 1560 -160 1650 -150
rect 1560 -730 1570 -160
rect 1590 -730 1620 -160
rect 1640 -730 1650 -160
rect 1560 -740 1650 -730
rect 60 -800 1500 -760
<< viali >>
rect -80 1455 -60 2025
rect -30 1455 -10 2025
rect 170 1455 190 2025
rect 1370 1455 1390 2025
rect 770 1385 790 1405
rect 1015 1385 1045 1405
rect 1570 1455 1590 2025
rect 1620 1455 1640 2025
rect 40 1345 90 1365
rect 1470 1345 1520 1365
rect -80 730 -60 1300
rect -30 730 -10 1300
rect 670 730 690 1300
rect 770 730 790 1300
rect 870 730 890 1300
rect 120 670 140 690
rect 520 670 540 690
rect 1420 670 1440 690
rect 1570 730 1590 1300
rect 1620 730 1640 1300
rect -80 -5 -60 565
rect -30 -5 -10 565
rect 120 605 140 625
rect 1020 605 1040 625
rect 1420 605 1440 625
rect 670 -5 690 565
rect 770 -5 790 565
rect 870 -5 890 565
rect 1570 -5 1590 565
rect 1620 -5 1640 565
rect -80 -730 -60 -160
rect -30 -730 -10 -160
rect 215 -110 245 -90
rect 515 -110 545 -90
rect 1315 -110 1345 -90
rect 170 -730 190 -160
rect 1370 -730 1390 -160
rect 1570 -730 1590 -160
rect 1620 -730 1640 -160
<< metal1 >>
rect -100 2025 1655 2035
rect -100 1455 -80 2025
rect -60 1455 -30 2025
rect -10 1455 170 2025
rect 190 1455 1370 2025
rect 1390 1455 1570 2025
rect 1590 1455 1620 2025
rect 1640 1455 1655 2025
rect -100 1445 1655 1455
rect -95 1300 0 1445
rect -95 730 -80 1300
rect -60 730 -30 1300
rect -10 730 0 1300
rect -95 720 0 730
rect 30 1365 100 1375
rect 30 1345 40 1365
rect 90 1345 100 1365
rect 30 1335 100 1345
rect 30 635 70 1335
rect 605 1300 700 1445
rect 605 730 670 1300
rect 690 730 700 1300
rect 605 720 700 730
rect 760 1405 800 1415
rect 760 1385 770 1405
rect 790 1385 800 1405
rect 760 1300 800 1385
rect 760 730 770 1300
rect 790 730 800 1300
rect 105 690 255 700
rect 105 670 120 690
rect 140 670 255 690
rect 105 660 255 670
rect 30 625 155 635
rect 30 605 120 625
rect 140 605 155 625
rect 30 595 155 605
rect -95 565 0 575
rect -95 -5 -80 565
rect -60 -5 -30 565
rect -10 -5 0 565
rect -95 -150 0 -5
rect 205 -90 255 660
rect 205 -110 215 -90
rect 245 -110 255 -90
rect 205 -120 255 -110
rect 505 690 555 700
rect 505 670 520 690
rect 540 670 555 690
rect 505 -90 555 670
rect 505 -110 515 -90
rect 545 -110 555 -90
rect 505 -120 555 -110
rect 605 565 700 575
rect 605 -5 670 565
rect 690 -5 700 565
rect 605 -150 700 -5
rect 760 565 800 730
rect 860 1300 955 1445
rect 860 730 870 1300
rect 890 730 955 1300
rect 860 720 955 730
rect 1005 1405 1055 1415
rect 1005 1385 1015 1405
rect 1045 1385 1055 1405
rect 1005 625 1055 1385
rect 1460 1365 1530 1375
rect 1460 1345 1470 1365
rect 1520 1345 1530 1365
rect 1460 1335 1530 1345
rect 1005 605 1020 625
rect 1040 605 1055 625
rect 1005 595 1055 605
rect 1305 690 1455 700
rect 1305 670 1420 690
rect 1440 670 1455 690
rect 1305 660 1455 670
rect 760 -5 770 565
rect 790 -5 800 565
rect 760 -15 800 -5
rect 860 565 955 575
rect 860 -5 870 565
rect 890 -5 955 565
rect 860 -150 955 -5
rect 1305 -90 1355 660
rect 1490 635 1530 1335
rect 1560 1300 1655 1445
rect 1560 730 1570 1300
rect 1590 730 1620 1300
rect 1640 730 1655 1300
rect 1560 720 1655 730
rect 1405 625 1530 635
rect 1405 605 1420 625
rect 1440 605 1530 625
rect 1405 595 1530 605
rect 1305 -110 1315 -90
rect 1345 -110 1355 -90
rect 1305 -120 1355 -110
rect 1560 565 1655 575
rect 1560 -5 1570 565
rect 1590 -5 1620 565
rect 1640 -5 1655 565
rect 1560 -150 1655 -5
rect -95 -160 1655 -150
rect -95 -730 -80 -160
rect -60 -730 -30 -160
rect -10 -730 170 -160
rect 190 -730 1370 -160
rect 1390 -730 1570 -160
rect 1590 -730 1620 -160
rect 1640 -730 1655 -160
rect -95 -740 1655 -730
<< labels >>
rlabel poly 1655 2085 1655 2085 3 Vbp
port 1 e
rlabel metal1 1655 1740 1655 1740 3 VP
port 2 e
rlabel poly 1655 1345 1655 1345 3 Vcp
port 3 e
rlabel poly 1655 -50 1655 -50 3 Vcn
port 4 e
rlabel metal1 1655 -445 1655 -445 3 VN
port 5 e
rlabel poly 1655 -790 1655 -790 3 Vbn
port 6 e
<< end >>
