magic
tech sky130A
timestamp 1697134827
<< nwell >>
rect -120 1245 1020 1885
<< nmos >>
rect 0 530 50 1130
rect 100 530 150 1130
rect 200 530 250 1130
rect 300 530 350 1130
rect 400 530 450 1130
rect 500 530 550 1130
rect 600 530 650 1130
rect 700 530 750 1130
rect 800 530 850 1130
rect 900 530 950 1130
rect 0 95 50 395
rect 100 95 150 395
rect 200 95 250 395
rect 300 95 350 395
rect 400 95 450 395
rect 500 95 550 395
rect 600 95 650 395
rect 700 95 750 395
rect 800 95 850 395
rect 900 95 950 395
rect 0 -310 50 -10
rect 100 -310 150 -10
rect 200 -310 250 -10
rect 300 -310 350 -10
rect 400 -310 450 -10
rect 500 -310 550 -10
rect 600 -310 650 -10
rect 700 -310 750 -10
rect 800 -310 850 -10
rect 900 -310 950 -10
<< pmos >>
rect 0 1265 50 1865
rect 100 1265 150 1865
rect 200 1265 250 1865
rect 300 1265 350 1865
rect 400 1265 450 1865
rect 500 1265 550 1865
rect 600 1265 650 1865
rect 700 1265 750 1865
rect 800 1265 850 1865
rect 900 1265 950 1865
<< ndiff >>
rect -50 1115 0 1130
rect -50 545 -35 1115
rect -15 545 0 1115
rect -50 530 0 545
rect 50 1115 100 1130
rect 50 545 65 1115
rect 85 545 100 1115
rect 50 530 100 545
rect 150 530 200 1130
rect 250 1115 300 1130
rect 250 545 265 1115
rect 285 545 300 1115
rect 250 530 300 545
rect 350 530 400 1130
rect 450 1115 500 1130
rect 450 545 465 1115
rect 485 545 500 1115
rect 450 530 500 545
rect 550 530 600 1130
rect 650 1115 700 1130
rect 650 545 665 1115
rect 685 545 700 1115
rect 650 530 700 545
rect 750 530 800 1130
rect 850 1115 900 1130
rect 850 545 865 1115
rect 885 545 900 1115
rect 850 530 900 545
rect 950 1115 1000 1130
rect 950 545 965 1115
rect 985 545 1000 1115
rect 950 530 1000 545
rect -50 380 0 395
rect -50 110 -35 380
rect -15 110 0 380
rect -50 95 0 110
rect 50 380 100 395
rect 50 110 65 380
rect 85 110 100 380
rect 50 95 100 110
rect 150 380 200 395
rect 150 110 165 380
rect 185 110 200 380
rect 150 95 200 110
rect 250 380 300 395
rect 250 110 265 380
rect 285 110 300 380
rect 250 95 300 110
rect 350 380 400 395
rect 350 110 365 380
rect 385 110 400 380
rect 350 95 400 110
rect 450 380 500 395
rect 450 110 465 380
rect 485 110 500 380
rect 450 95 500 110
rect 550 380 600 395
rect 550 110 565 380
rect 585 110 600 380
rect 550 95 600 110
rect 650 380 700 395
rect 650 110 665 380
rect 685 110 700 380
rect 650 95 700 110
rect 750 380 800 395
rect 750 110 765 380
rect 785 110 800 380
rect 750 95 800 110
rect 850 380 900 395
rect 850 110 865 380
rect 885 110 900 380
rect 850 95 900 110
rect 950 380 1000 395
rect 950 110 965 380
rect 985 110 1000 380
rect 950 95 1000 110
rect -50 -25 0 -10
rect -50 -295 -35 -25
rect -15 -295 0 -25
rect -50 -310 0 -295
rect 50 -25 100 -10
rect 50 -295 65 -25
rect 85 -295 100 -25
rect 50 -310 100 -295
rect 150 -25 200 -10
rect 150 -295 165 -25
rect 185 -295 200 -25
rect 150 -310 200 -295
rect 250 -25 300 -10
rect 250 -295 265 -25
rect 285 -295 300 -25
rect 250 -310 300 -295
rect 350 -25 400 -10
rect 350 -295 365 -25
rect 385 -295 400 -25
rect 350 -310 400 -295
rect 450 -25 500 -10
rect 450 -295 465 -25
rect 485 -295 500 -25
rect 450 -310 500 -295
rect 550 -25 600 -10
rect 550 -295 565 -25
rect 585 -295 600 -25
rect 550 -310 600 -295
rect 650 -25 700 -10
rect 650 -295 665 -25
rect 685 -295 700 -25
rect 650 -310 700 -295
rect 750 -25 800 -10
rect 750 -295 765 -25
rect 785 -295 800 -25
rect 750 -310 800 -295
rect 850 -25 900 -10
rect 850 -295 865 -25
rect 885 -295 900 -25
rect 850 -310 900 -295
rect 950 -25 1000 -10
rect 950 -295 965 -25
rect 985 -295 1000 -25
rect 950 -310 1000 -295
<< pdiff >>
rect -50 1850 0 1865
rect -50 1280 -35 1850
rect -15 1280 0 1850
rect -50 1265 0 1280
rect 50 1850 100 1865
rect 50 1280 65 1850
rect 85 1280 100 1850
rect 50 1265 100 1280
rect 150 1850 200 1865
rect 150 1280 165 1850
rect 185 1280 200 1850
rect 150 1265 200 1280
rect 250 1850 300 1865
rect 250 1280 265 1850
rect 285 1280 300 1850
rect 250 1265 300 1280
rect 350 1850 400 1865
rect 350 1280 365 1850
rect 385 1280 400 1850
rect 350 1265 400 1280
rect 450 1850 500 1865
rect 450 1280 465 1850
rect 485 1280 500 1850
rect 450 1265 500 1280
rect 550 1850 600 1865
rect 550 1280 565 1850
rect 585 1280 600 1850
rect 550 1265 600 1280
rect 650 1850 700 1865
rect 650 1280 665 1850
rect 685 1280 700 1850
rect 650 1265 700 1280
rect 750 1850 800 1865
rect 750 1280 765 1850
rect 785 1280 800 1850
rect 750 1265 800 1280
rect 850 1850 900 1865
rect 850 1280 865 1850
rect 885 1280 900 1850
rect 850 1265 900 1280
rect 950 1850 1000 1865
rect 950 1280 965 1850
rect 985 1280 1000 1850
rect 950 1265 1000 1280
<< ndiffc >>
rect -35 545 -15 1115
rect 65 545 85 1115
rect 265 545 285 1115
rect 465 545 485 1115
rect 665 545 685 1115
rect 865 545 885 1115
rect 965 545 985 1115
rect -35 110 -15 380
rect 65 110 85 380
rect 165 110 185 380
rect 265 110 285 380
rect 365 110 385 380
rect 465 110 485 380
rect 565 110 585 380
rect 665 110 685 380
rect 765 110 785 380
rect 865 110 885 380
rect 965 110 985 380
rect -35 -295 -15 -25
rect 65 -295 85 -25
rect 165 -295 185 -25
rect 265 -295 285 -25
rect 365 -295 385 -25
rect 465 -295 485 -25
rect 565 -295 585 -25
rect 665 -295 685 -25
rect 765 -295 785 -25
rect 865 -295 885 -25
rect 965 -295 985 -25
<< pdiffc >>
rect -35 1280 -15 1850
rect 65 1280 85 1850
rect 165 1280 185 1850
rect 265 1280 285 1850
rect 365 1280 385 1850
rect 465 1280 485 1850
rect 565 1280 585 1850
rect 665 1280 685 1850
rect 765 1280 785 1850
rect 865 1280 885 1850
rect 965 1280 985 1850
<< psubdiff >>
rect -100 1115 -50 1130
rect -100 545 -85 1115
rect -65 545 -50 1115
rect -100 530 -50 545
rect -100 380 -50 395
rect -100 110 -85 380
rect -65 110 -50 380
rect -100 95 -50 110
rect -100 -25 -50 -10
rect -100 -295 -85 -25
rect -65 -295 -50 -25
rect -100 -310 -50 -295
<< nsubdiff >>
rect -100 1850 -50 1865
rect -100 1280 -85 1850
rect -65 1280 -50 1850
rect -100 1265 -50 1280
<< psubdiffcont >>
rect -85 545 -65 1115
rect -85 110 -65 380
rect -85 -295 -65 -25
<< nsubdiffcont >>
rect -85 1280 -65 1850
<< poly >>
rect -95 1905 750 1920
rect 0 1865 50 1880
rect 100 1865 150 1880
rect 200 1865 250 1905
rect 300 1865 350 1905
rect 400 1865 450 1880
rect 500 1865 550 1880
rect 600 1865 650 1905
rect 700 1865 750 1905
rect 800 1865 850 1880
rect 900 1865 950 1880
rect 0 1250 50 1265
rect -95 1240 50 1250
rect -95 1220 -85 1240
rect -65 1235 50 1240
rect -65 1220 -55 1235
rect 100 1225 150 1265
rect 200 1250 250 1265
rect 300 1250 350 1265
rect 400 1225 450 1265
rect 500 1225 550 1265
rect 600 1250 650 1265
rect 700 1250 750 1265
rect 800 1225 850 1265
rect 900 1250 950 1265
rect 900 1240 995 1250
rect 900 1235 965 1240
rect -95 1210 -55 1220
rect 75 1210 850 1225
rect 955 1220 965 1235
rect 985 1220 995 1240
rect 955 1210 995 1220
rect 75 1205 90 1210
rect 30 1190 90 1205
rect 30 1185 45 1190
rect -100 1170 45 1185
rect 120 1170 850 1185
rect 0 1130 50 1145
rect 100 1130 150 1170
rect 200 1130 250 1145
rect 300 1130 350 1145
rect 400 1130 450 1170
rect 500 1130 550 1170
rect 600 1130 650 1145
rect 700 1130 750 1145
rect 800 1130 850 1170
rect 955 1175 995 1185
rect 955 1160 965 1175
rect 900 1155 965 1160
rect 985 1155 995 1175
rect 900 1145 995 1155
rect 900 1130 950 1145
rect 0 515 50 530
rect -95 505 50 515
rect -95 485 -85 505
rect -65 500 50 505
rect -65 485 -55 500
rect 100 490 150 530
rect -95 475 -55 485
rect 75 475 150 490
rect 200 505 250 530
rect 200 485 215 505
rect 235 485 250 505
rect 200 475 250 485
rect 300 505 350 530
rect 400 515 450 530
rect 500 515 550 530
rect 300 485 315 505
rect 335 485 350 505
rect 300 475 350 485
rect 600 505 650 530
rect 600 485 615 505
rect 635 485 650 505
rect 600 475 650 485
rect 700 505 750 530
rect 800 515 850 530
rect 900 515 950 530
rect 700 485 715 505
rect 735 485 750 505
rect 700 475 750 485
rect 860 475 1000 490
rect 30 460 90 475
rect 30 450 45 460
rect 860 450 875 475
rect -100 435 45 450
rect 120 435 875 450
rect 955 440 995 450
rect 0 395 50 410
rect 100 395 150 435
rect 200 395 250 410
rect 300 395 350 410
rect 400 395 450 435
rect 500 395 550 435
rect 600 395 650 410
rect 700 395 750 410
rect 800 395 850 435
rect 955 425 965 440
rect 900 420 965 425
rect 985 420 995 440
rect 900 410 995 420
rect 900 395 950 410
rect 0 80 50 95
rect 100 80 150 95
rect -95 70 50 80
rect -95 50 -85 70
rect -65 65 50 70
rect -65 50 -55 65
rect -95 40 -55 50
rect 200 55 250 95
rect 300 55 350 95
rect 400 80 450 95
rect 500 80 550 95
rect 600 55 650 95
rect 700 55 750 95
rect 800 80 850 95
rect 900 80 950 95
rect 200 40 1000 55
rect 0 30 50 40
rect 0 10 10 30
rect 30 10 50 30
rect 0 -10 50 10
rect 100 -10 150 5
rect 200 -10 250 5
rect 300 -10 350 5
rect 400 -10 450 5
rect 500 -10 550 5
rect 600 -10 650 5
rect 700 -10 750 5
rect 800 -10 850 5
rect 900 -10 950 5
rect 0 -325 50 -310
rect 100 -335 150 -310
rect 100 -355 115 -335
rect 135 -355 150 -335
rect 100 -365 150 -355
rect 200 -335 250 -310
rect 200 -355 215 -335
rect 235 -355 250 -335
rect 200 -365 250 -355
rect 300 -335 350 -310
rect 300 -355 315 -335
rect 335 -355 350 -335
rect 300 -365 350 -355
rect 400 -335 450 -310
rect 400 -355 415 -335
rect 435 -355 450 -335
rect 400 -365 450 -355
rect 500 -335 550 -310
rect 500 -355 515 -335
rect 535 -355 550 -335
rect 500 -365 550 -355
rect 600 -335 650 -310
rect 600 -355 615 -335
rect 635 -355 650 -335
rect 600 -365 650 -355
rect 700 -335 750 -310
rect 700 -355 715 -335
rect 735 -355 750 -335
rect 700 -365 750 -355
rect 800 -335 850 -310
rect 800 -355 815 -335
rect 835 -355 850 -335
rect 900 -325 950 -310
rect 900 -335 995 -325
rect 900 -340 965 -335
rect 800 -365 850 -355
rect 955 -355 965 -340
rect 985 -355 995 -335
rect 955 -365 995 -355
<< polycont >>
rect -85 1220 -65 1240
rect 965 1220 985 1240
rect 965 1155 985 1175
rect -85 485 -65 505
rect 215 485 235 505
rect 315 485 335 505
rect 615 485 635 505
rect 715 485 735 505
rect 965 420 985 440
rect -85 50 -65 70
rect 10 10 30 30
rect 115 -355 135 -335
rect 215 -355 235 -335
rect 315 -355 335 -335
rect 415 -355 435 -335
rect 515 -355 535 -335
rect 615 -355 635 -335
rect 715 -355 735 -335
rect 815 -355 835 -335
rect 965 -355 985 -335
<< locali >>
rect 455 1880 1000 1920
rect -95 1850 -5 1860
rect -95 1280 -85 1850
rect -65 1280 -35 1850
rect -15 1280 -5 1850
rect -95 1270 -5 1280
rect 55 1850 95 1860
rect 55 1280 65 1850
rect 85 1280 95 1850
rect -95 1240 -55 1270
rect -95 1220 -85 1240
rect -65 1220 -55 1240
rect -95 1210 -55 1220
rect -95 1115 -5 1125
rect -95 545 -85 1115
rect -65 545 -35 1115
rect -15 545 -5 1115
rect -95 535 -5 545
rect 55 1115 95 1280
rect 55 545 65 1115
rect 85 545 95 1115
rect -95 505 -55 535
rect -95 485 -85 505
rect -65 485 -55 505
rect -95 475 -55 485
rect 55 515 95 545
rect 155 1850 195 1860
rect 155 1280 165 1850
rect 185 1280 195 1850
rect 155 585 195 1280
rect 255 1850 295 1860
rect 255 1280 265 1850
rect 285 1280 295 1850
rect 255 1270 295 1280
rect 355 1850 395 1860
rect 355 1280 365 1850
rect 385 1280 395 1850
rect 155 545 165 585
rect 185 545 195 585
rect 155 535 195 545
rect 255 1115 295 1125
rect 255 545 265 1115
rect 285 545 295 1115
rect 255 535 295 545
rect 355 585 395 1280
rect 355 545 365 585
rect 385 545 395 585
rect 355 535 395 545
rect 455 1850 495 1880
rect 455 1280 465 1850
rect 485 1280 495 1850
rect 455 1115 495 1280
rect 455 545 465 1115
rect 485 545 495 1115
rect 455 535 495 545
rect 555 1850 595 1860
rect 555 1280 565 1850
rect 585 1280 595 1850
rect 555 585 595 1280
rect 655 1850 695 1860
rect 655 1280 665 1850
rect 685 1280 695 1850
rect 655 1270 695 1280
rect 755 1850 795 1860
rect 755 1280 765 1850
rect 785 1280 795 1850
rect 555 545 565 585
rect 585 545 595 585
rect 555 535 595 545
rect 655 1115 695 1125
rect 655 545 665 1115
rect 685 545 695 1115
rect 655 535 695 545
rect 755 585 795 1280
rect 755 545 765 585
rect 785 545 795 585
rect 755 535 795 545
rect 855 1850 895 1860
rect 855 1280 865 1850
rect 885 1280 895 1850
rect 855 1115 895 1280
rect 955 1850 1000 1860
rect 955 1280 965 1850
rect 985 1280 1000 1850
rect 955 1270 1000 1280
rect 955 1240 995 1270
rect 955 1220 965 1240
rect 985 1220 995 1240
rect 955 1210 995 1220
rect 855 545 865 1115
rect 885 545 895 1115
rect 855 515 895 545
rect 955 1175 995 1185
rect 955 1155 965 1175
rect 985 1155 995 1175
rect 955 1125 995 1155
rect 955 1115 1000 1125
rect 955 545 965 1115
rect 985 545 1000 1115
rect 955 535 1000 545
rect 55 505 895 515
rect 55 485 215 505
rect 235 485 315 505
rect 335 485 615 505
rect 635 485 715 505
rect 735 485 895 505
rect 55 475 895 485
rect 55 440 895 450
rect 55 420 155 440
rect 195 420 755 440
rect 795 420 895 440
rect 55 410 895 420
rect -95 380 -5 390
rect -95 110 -85 380
rect -65 110 -35 380
rect -15 110 -5 380
rect -95 100 -5 110
rect 55 380 95 410
rect 55 110 65 380
rect 85 110 95 380
rect 55 100 95 110
rect 155 380 195 390
rect 155 110 165 380
rect 185 110 195 380
rect -95 70 -55 100
rect -95 50 -85 70
rect -65 50 -55 70
rect -95 40 -55 50
rect 155 70 195 110
rect 255 380 295 390
rect 255 110 265 380
rect 285 110 295 380
rect 255 100 295 110
rect 355 380 395 390
rect 355 110 365 380
rect 385 110 395 380
rect 355 70 395 110
rect 455 380 495 410
rect 455 110 465 380
rect 485 110 495 380
rect 455 100 495 110
rect 555 380 595 390
rect 555 110 565 380
rect 585 110 595 380
rect 555 70 595 110
rect 655 380 695 390
rect 655 110 665 380
rect 685 110 695 380
rect 655 100 695 110
rect 755 380 795 390
rect 755 110 765 380
rect 785 110 795 380
rect 755 70 795 110
rect 855 380 895 410
rect 855 110 865 380
rect 885 110 895 380
rect 855 100 895 110
rect 955 440 995 450
rect 955 420 965 440
rect 985 420 995 440
rect 955 390 995 420
rect 955 380 1000 390
rect 955 110 965 380
rect 985 110 1000 380
rect 955 100 1000 110
rect -35 30 40 40
rect 155 30 795 70
rect -35 10 10 30
rect 30 10 40 30
rect -35 0 40 10
rect -35 -15 -5 0
rect -95 -25 -5 -15
rect -95 -295 -85 -25
rect -65 -295 -35 -25
rect -15 -295 -5 -25
rect -95 -305 -5 -295
rect 55 -25 95 -15
rect 55 -295 65 -25
rect 85 -295 95 -25
rect 55 -325 95 -295
rect 155 -25 195 -15
rect 155 -295 165 -25
rect 185 -295 195 -25
rect 155 -305 195 -295
rect 255 -25 295 30
rect 255 -295 265 -25
rect 285 -295 295 -25
rect 255 -305 295 -295
rect 355 -25 395 -15
rect 355 -295 365 -25
rect 385 -295 395 -25
rect 355 -305 395 -295
rect 455 -25 495 -15
rect 455 -295 465 -25
rect 485 -295 495 -25
rect 455 -325 495 -295
rect 555 -25 595 -15
rect 555 -295 565 -25
rect 585 -295 595 -25
rect 555 -305 595 -295
rect 655 -25 695 30
rect 655 -295 665 -25
rect 685 -295 695 -25
rect 655 -305 695 -295
rect 755 -25 795 -15
rect 755 -295 765 -25
rect 785 -295 795 -25
rect 755 -305 795 -295
rect 855 -25 895 -15
rect 855 -295 865 -25
rect 885 -295 895 -25
rect 855 -325 895 -295
rect -100 -335 895 -325
rect -100 -355 115 -335
rect 135 -355 215 -335
rect 235 -355 315 -335
rect 335 -355 415 -335
rect 435 -355 515 -335
rect 535 -355 615 -335
rect 635 -355 715 -335
rect 735 -355 815 -335
rect 835 -355 895 -335
rect -100 -365 895 -355
rect 955 -25 1000 -15
rect 955 -295 965 -25
rect 985 -295 1000 -25
rect 955 -305 1000 -295
rect 955 -335 995 -305
rect 955 -355 965 -335
rect 985 -355 995 -335
rect 955 -365 995 -355
<< viali >>
rect -85 1280 -65 1850
rect -35 1280 -15 1850
rect -85 545 -65 1115
rect -35 545 -15 1115
rect 265 1280 285 1850
rect 165 545 185 585
rect 265 545 285 1115
rect 365 545 385 585
rect 665 1280 685 1850
rect 565 545 585 585
rect 665 545 685 1115
rect 765 545 785 585
rect 965 1280 985 1850
rect 965 545 985 1115
rect 155 420 195 440
rect 755 420 795 440
rect -85 110 -65 380
rect -35 110 -15 380
rect 265 110 285 380
rect 665 110 685 380
rect 965 110 985 380
rect -85 -295 -65 -25
rect -35 -295 -15 -25
rect 165 -295 185 -25
rect 365 -295 385 -25
rect 565 -295 585 -25
rect 765 -295 785 -25
rect 965 -295 985 -25
<< metal1 >>
rect -100 1850 1000 1860
rect -100 1280 -85 1850
rect -65 1280 -35 1850
rect -15 1280 265 1850
rect 285 1280 665 1850
rect 685 1280 965 1850
rect 985 1280 1000 1850
rect -100 1270 1000 1280
rect -100 1115 1000 1125
rect -100 545 -85 1115
rect -65 545 -35 1115
rect -15 625 265 1115
rect -15 545 125 625
rect -100 535 125 545
rect 155 585 195 595
rect 155 545 165 585
rect 185 545 195 585
rect -100 380 -5 535
rect 155 450 195 545
rect 225 545 265 625
rect 285 625 665 1115
rect 285 545 325 625
rect 225 535 325 545
rect 355 585 395 595
rect 355 545 365 585
rect 385 545 395 585
rect 145 440 205 450
rect 145 420 155 440
rect 195 420 205 440
rect 145 410 205 420
rect 355 390 395 545
rect 555 585 595 595
rect 555 545 565 585
rect 585 545 595 585
rect 555 390 595 545
rect 625 545 665 625
rect 685 625 965 1115
rect 685 545 725 625
rect 625 535 725 545
rect 755 585 795 595
rect 755 545 765 585
rect 785 545 795 585
rect 755 450 795 545
rect 825 545 965 625
rect 985 545 1000 1115
rect 825 535 1000 545
rect 745 440 805 450
rect 745 420 755 440
rect 795 420 805 440
rect 745 410 805 420
rect -100 110 -85 380
rect -65 110 -35 380
rect -15 110 -5 380
rect -100 -15 -5 110
rect 255 380 900 390
rect 255 110 265 380
rect 285 110 665 380
rect 685 110 900 380
rect 255 100 900 110
rect 955 380 1000 535
rect 955 110 965 380
rect 985 110 1000 380
rect 955 -15 1000 110
rect -100 -25 1000 -15
rect -100 -295 -85 -25
rect -65 -295 -35 -25
rect -15 -295 165 -25
rect 185 -295 365 -25
rect 385 -295 565 -25
rect 585 -295 765 -25
rect 785 -295 965 -25
rect 985 -295 1000 -25
rect -100 -305 1000 -295
<< labels >>
rlabel poly -100 445 -100 445 7 Vcn
port 2 w
rlabel locali -100 -345 -100 -345 7 Vbn
port 1 w
rlabel metal1 -100 980 -100 980 7 VN
port 3 w
rlabel poly -100 1175 -100 1175 7 Vcp
port 4 w
rlabel metal1 -100 1715 -100 1715 7 VP
port 5 w
rlabel poly -95 1910 -95 1910 7 Vbp
port 6 w
rlabel locali 1000 1900 1000 1900 3 Vout
port 7 e
rlabel poly 1000 485 1000 485 3 V1
port 8 e
rlabel poly 1000 45 1000 45 3 V2
port 9 e
<< end >>
