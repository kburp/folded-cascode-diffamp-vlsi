magic
tech sky130A
timestamp 1697131150
<< poly >>
rect 1770 2880 1810 2895
rect 1795 2195 1810 2880
rect 1795 2180 1840 2195
rect 1770 2140 1800 2155
rect 1785 950 1800 2140
rect 1825 1385 1840 2180
rect 1825 1370 1850 1385
rect 1785 935 1830 950
rect 1770 740 1810 755
rect 1795 515 1810 740
rect 1795 500 1840 515
rect 1830 30 1870 40
rect 1830 15 1840 30
rect 1770 10 1840 15
rect 1860 10 1870 30
rect 1770 0 1870 10
<< polycont >>
rect 1840 10 1860 30
<< metal1 >>
rect 1720 1465 1770 1520
rect 1720 1415 1880 1465
rect 1830 1325 1880 1415
rect 1770 60 1830 890
use biasgen  biasgen_0
timestamp 1697129952
transform 1 0 115 0 1 800
box -115 -800 1675 2095
use fc_diffamp  fc_diffamp_0
timestamp 1697130813
transform 1 0 1930 0 1 65
box -120 -65 1870 1320
<< end >>
