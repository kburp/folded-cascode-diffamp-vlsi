magic
tech sky130A
timestamp 1697135791
<< nwell >>
rect 1790 2155 1800 2250
rect 1770 2140 1800 2155
rect 1790 1610 1800 2140
<< poly >>
rect 1770 2880 1800 2895
rect 1780 2285 1800 2880
rect 1780 2270 1825 2285
rect 1770 2140 1795 2155
rect 1780 1550 1795 2140
rect 1780 1535 1825 1550
rect 1780 800 1815 815
rect 1780 755 1795 800
rect 1770 740 1795 755
rect 1815 30 1855 40
rect 1815 15 1825 30
rect 1770 10 1825 15
rect 1845 10 1855 30
rect 1770 0 1855 10
<< polycont >>
rect 1825 10 1845 30
<< metal1 >>
rect 1765 1635 1815 2225
rect 1770 60 1815 1375
use biasgen  biasgen_0
timestamp 1697129952
transform 1 0 115 0 1 800
box -115 -800 1675 2095
use fc_diffamp  fc_diffamp_0
timestamp 1697134827
transform 1 0 1915 0 1 365
box -120 -365 1020 1920
<< labels >>
rlabel space 2915 2265 2915 2265 3 Vout
rlabel space 2915 850 2915 850 3 V1
rlabel space 2915 410 2915 410 3 V2
rlabel space 2915 210 2915 210 1 VN
rlabel space 2915 1930 2915 1930 1 VP
<< end >>
