magic
tech sky130A
timestamp 1697129871
<< nwell >>
rect -120 945 1870 1285
<< nmos >>
rect 0 530 50 830
rect 100 530 150 830
rect 200 530 250 830
rect 300 530 350 830
rect 400 530 450 830
rect 500 530 550 830
rect 600 530 650 830
rect 700 530 750 830
rect 800 530 850 830
rect 900 530 950 830
rect 1000 530 1050 830
rect 1100 530 1150 830
rect 1200 530 1250 830
rect 1300 530 1350 830
rect 1400 530 1450 830
rect 1500 530 1550 830
rect 1600 530 1650 830
rect 1700 530 1750 830
rect 0 245 50 395
rect 100 245 150 395
rect 200 245 250 395
rect 300 245 350 395
rect 400 245 450 395
rect 500 245 550 395
rect 600 245 650 395
rect 700 245 750 395
rect 800 245 850 395
rect 900 245 950 395
rect 1000 245 1050 395
rect 1100 245 1150 395
rect 1200 245 1250 395
rect 1300 245 1350 395
rect 1400 245 1450 395
rect 1500 245 1550 395
rect 1600 245 1650 395
rect 1700 245 1750 395
rect 0 -10 50 140
rect 100 -10 150 140
rect 200 -10 250 140
rect 300 -10 350 140
rect 400 -10 450 140
rect 500 -10 550 140
rect 600 -10 650 140
rect 700 -10 750 140
rect 800 -10 850 140
rect 900 -10 950 140
rect 1000 -10 1050 140
rect 1100 -10 1150 140
rect 1200 -10 1250 140
rect 1300 -10 1350 140
rect 1400 -10 1450 140
rect 1500 -10 1550 140
rect 1600 -10 1650 140
rect 1700 -10 1750 140
<< pmos >>
rect 0 965 50 1265
rect 100 965 150 1265
rect 200 965 250 1265
rect 300 965 350 1265
rect 400 965 450 1265
rect 500 965 550 1265
rect 600 965 650 1265
rect 700 965 750 1265
rect 800 965 850 1265
rect 900 965 950 1265
rect 1000 965 1050 1265
rect 1100 965 1150 1265
rect 1200 965 1250 1265
rect 1300 965 1350 1265
rect 1400 965 1450 1265
rect 1500 965 1550 1265
rect 1600 965 1650 1265
rect 1700 965 1750 1265
<< ndiff >>
rect -50 815 0 830
rect -50 545 -35 815
rect -15 545 0 815
rect -50 530 0 545
rect 50 815 100 830
rect 50 545 65 815
rect 85 545 100 815
rect 50 530 100 545
rect 150 530 200 830
rect 250 815 300 830
rect 250 545 265 815
rect 285 545 300 815
rect 250 530 300 545
rect 350 530 400 830
rect 450 815 500 830
rect 450 545 465 815
rect 485 545 500 815
rect 450 530 500 545
rect 550 530 600 830
rect 650 815 700 830
rect 650 545 665 815
rect 685 545 700 815
rect 650 530 700 545
rect 750 530 800 830
rect 850 815 900 830
rect 850 545 865 815
rect 885 545 900 815
rect 850 530 900 545
rect 950 530 1000 830
rect 1050 815 1100 830
rect 1050 545 1065 815
rect 1085 545 1100 815
rect 1050 530 1100 545
rect 1150 530 1200 830
rect 1250 815 1300 830
rect 1250 545 1265 815
rect 1285 545 1300 815
rect 1250 530 1300 545
rect 1350 530 1400 830
rect 1450 815 1500 830
rect 1450 545 1465 815
rect 1485 545 1500 815
rect 1450 530 1500 545
rect 1550 530 1600 830
rect 1650 815 1700 830
rect 1650 545 1665 815
rect 1685 545 1700 815
rect 1650 530 1700 545
rect 1750 815 1800 830
rect 1750 545 1765 815
rect 1785 545 1800 815
rect 1750 530 1800 545
rect -50 380 0 395
rect -50 260 -35 380
rect -15 260 0 380
rect -50 245 0 260
rect 50 380 100 395
rect 50 260 65 380
rect 85 260 100 380
rect 50 245 100 260
rect 150 380 200 395
rect 150 260 165 380
rect 185 260 200 380
rect 150 245 200 260
rect 250 380 300 395
rect 250 260 265 380
rect 285 260 300 380
rect 250 245 300 260
rect 350 380 400 395
rect 350 260 365 380
rect 385 260 400 380
rect 350 245 400 260
rect 450 380 500 395
rect 450 260 465 380
rect 485 260 500 380
rect 450 245 500 260
rect 550 380 600 395
rect 550 260 565 380
rect 585 260 600 380
rect 550 245 600 260
rect 650 380 700 395
rect 650 260 665 380
rect 685 260 700 380
rect 650 245 700 260
rect 750 380 800 395
rect 750 260 765 380
rect 785 260 800 380
rect 750 245 800 260
rect 850 380 900 395
rect 850 260 865 380
rect 885 260 900 380
rect 850 245 900 260
rect 950 380 1000 395
rect 950 260 965 380
rect 985 260 1000 380
rect 950 245 1000 260
rect 1050 380 1100 395
rect 1050 260 1065 380
rect 1085 260 1100 380
rect 1050 245 1100 260
rect 1150 380 1200 395
rect 1150 260 1165 380
rect 1185 260 1200 380
rect 1150 245 1200 260
rect 1250 380 1300 395
rect 1250 260 1265 380
rect 1285 260 1300 380
rect 1250 245 1300 260
rect 1350 380 1400 395
rect 1350 260 1365 380
rect 1385 260 1400 380
rect 1350 245 1400 260
rect 1450 380 1500 395
rect 1450 260 1465 380
rect 1485 260 1500 380
rect 1450 245 1500 260
rect 1550 380 1600 395
rect 1550 260 1565 380
rect 1585 260 1600 380
rect 1550 245 1600 260
rect 1650 380 1700 395
rect 1650 260 1665 380
rect 1685 260 1700 380
rect 1650 245 1700 260
rect 1750 380 1800 395
rect 1750 260 1765 380
rect 1785 260 1800 380
rect 1750 245 1800 260
rect -50 125 0 140
rect -50 5 -35 125
rect -15 5 0 125
rect -50 -10 0 5
rect 50 125 100 140
rect 50 5 65 125
rect 85 5 100 125
rect 50 -10 100 5
rect 150 125 200 140
rect 150 5 165 125
rect 185 5 200 125
rect 150 -10 200 5
rect 250 125 300 140
rect 250 5 265 125
rect 285 5 300 125
rect 250 -10 300 5
rect 350 125 400 140
rect 350 5 365 125
rect 385 5 400 125
rect 350 -10 400 5
rect 450 125 500 140
rect 450 5 465 125
rect 485 5 500 125
rect 450 -10 500 5
rect 550 125 600 140
rect 550 5 565 125
rect 585 5 600 125
rect 550 -10 600 5
rect 650 125 700 140
rect 650 5 665 125
rect 685 5 700 125
rect 650 -10 700 5
rect 750 125 800 140
rect 750 5 765 125
rect 785 5 800 125
rect 750 -10 800 5
rect 850 125 900 140
rect 850 5 865 125
rect 885 5 900 125
rect 850 -10 900 5
rect 950 125 1000 140
rect 950 5 965 125
rect 985 5 1000 125
rect 950 -10 1000 5
rect 1050 125 1100 140
rect 1050 5 1065 125
rect 1085 5 1100 125
rect 1050 -10 1100 5
rect 1150 125 1200 140
rect 1150 5 1165 125
rect 1185 5 1200 125
rect 1150 -10 1200 5
rect 1250 125 1300 140
rect 1250 5 1265 125
rect 1285 5 1300 125
rect 1250 -10 1300 5
rect 1350 125 1400 140
rect 1350 5 1365 125
rect 1385 5 1400 125
rect 1350 -10 1400 5
rect 1450 125 1500 140
rect 1450 5 1465 125
rect 1485 5 1500 125
rect 1450 -10 1500 5
rect 1550 125 1600 140
rect 1550 5 1565 125
rect 1585 5 1600 125
rect 1550 -10 1600 5
rect 1650 125 1700 140
rect 1650 5 1665 125
rect 1685 5 1700 125
rect 1650 -10 1700 5
rect 1750 125 1800 140
rect 1750 5 1765 125
rect 1785 5 1800 125
rect 1750 -10 1800 5
<< pdiff >>
rect -50 1250 0 1265
rect -50 980 -35 1250
rect -15 980 0 1250
rect -50 965 0 980
rect 50 1250 100 1265
rect 50 980 65 1250
rect 85 980 100 1250
rect 50 965 100 980
rect 150 1250 200 1265
rect 150 980 165 1250
rect 185 980 200 1250
rect 150 965 200 980
rect 250 1250 300 1265
rect 250 980 265 1250
rect 285 980 300 1250
rect 250 965 300 980
rect 350 1250 400 1265
rect 350 980 365 1250
rect 385 980 400 1250
rect 350 965 400 980
rect 450 1250 500 1265
rect 450 980 465 1250
rect 485 980 500 1250
rect 450 965 500 980
rect 550 1250 600 1265
rect 550 980 565 1250
rect 585 980 600 1250
rect 550 965 600 980
rect 650 1250 700 1265
rect 650 980 665 1250
rect 685 980 700 1250
rect 650 965 700 980
rect 750 1250 800 1265
rect 750 980 765 1250
rect 785 980 800 1250
rect 750 965 800 980
rect 850 1250 900 1265
rect 850 980 865 1250
rect 885 980 900 1250
rect 850 965 900 980
rect 950 1250 1000 1265
rect 950 980 965 1250
rect 985 980 1000 1250
rect 950 965 1000 980
rect 1050 1250 1100 1265
rect 1050 980 1065 1250
rect 1085 980 1100 1250
rect 1050 965 1100 980
rect 1150 1250 1200 1265
rect 1150 980 1165 1250
rect 1185 980 1200 1250
rect 1150 965 1200 980
rect 1250 1250 1300 1265
rect 1250 980 1265 1250
rect 1285 980 1300 1250
rect 1250 965 1300 980
rect 1350 1250 1400 1265
rect 1350 980 1365 1250
rect 1385 980 1400 1250
rect 1350 965 1400 980
rect 1450 1250 1500 1265
rect 1450 980 1465 1250
rect 1485 980 1500 1250
rect 1450 965 1500 980
rect 1550 1250 1600 1265
rect 1550 980 1565 1250
rect 1585 980 1600 1250
rect 1550 965 1600 980
rect 1650 1250 1700 1265
rect 1650 980 1665 1250
rect 1685 980 1700 1250
rect 1650 965 1700 980
rect 1750 1250 1800 1265
rect 1750 980 1765 1250
rect 1785 980 1800 1250
rect 1750 965 1800 980
<< ndiffc >>
rect -35 545 -15 815
rect 65 545 85 815
rect 265 545 285 815
rect 465 545 485 815
rect 665 545 685 815
rect 865 545 885 815
rect 1065 545 1085 815
rect 1265 545 1285 815
rect 1465 545 1485 815
rect 1665 545 1685 815
rect 1765 545 1785 815
rect -35 260 -15 380
rect 65 260 85 380
rect 165 260 185 380
rect 265 260 285 380
rect 365 260 385 380
rect 465 260 485 380
rect 565 260 585 380
rect 665 260 685 380
rect 765 260 785 380
rect 865 260 885 380
rect 965 260 985 380
rect 1065 260 1085 380
rect 1165 260 1185 380
rect 1265 260 1285 380
rect 1365 260 1385 380
rect 1465 260 1485 380
rect 1565 260 1585 380
rect 1665 260 1685 380
rect 1765 260 1785 380
rect -35 5 -15 125
rect 65 5 85 125
rect 165 5 185 125
rect 265 5 285 125
rect 365 5 385 125
rect 465 5 485 125
rect 565 5 585 125
rect 665 5 685 125
rect 765 5 785 125
rect 865 5 885 125
rect 965 5 985 125
rect 1065 5 1085 125
rect 1165 5 1185 125
rect 1265 5 1285 125
rect 1365 5 1385 125
rect 1465 5 1485 125
rect 1565 5 1585 125
rect 1665 5 1685 125
rect 1765 5 1785 125
<< pdiffc >>
rect -35 980 -15 1250
rect 65 980 85 1250
rect 165 980 185 1250
rect 265 980 285 1250
rect 365 980 385 1250
rect 465 980 485 1250
rect 565 980 585 1250
rect 665 980 685 1250
rect 765 980 785 1250
rect 865 980 885 1250
rect 965 980 985 1250
rect 1065 980 1085 1250
rect 1165 980 1185 1250
rect 1265 980 1285 1250
rect 1365 980 1385 1250
rect 1465 980 1485 1250
rect 1565 980 1585 1250
rect 1665 980 1685 1250
rect 1765 980 1785 1250
<< psubdiff >>
rect -100 815 -50 830
rect -100 545 -85 815
rect -65 545 -50 815
rect -100 530 -50 545
rect 1800 815 1850 830
rect 1800 545 1815 815
rect 1835 545 1850 815
rect 1800 530 1850 545
rect -100 380 -50 395
rect -100 260 -85 380
rect -65 260 -50 380
rect -100 245 -50 260
rect 1800 380 1850 395
rect 1800 260 1815 380
rect 1835 260 1850 380
rect 1800 245 1850 260
rect -100 125 -50 140
rect -100 5 -85 125
rect -65 5 -50 125
rect -100 -10 -50 5
rect 1800 125 1850 140
rect 1800 5 1815 125
rect 1835 5 1850 125
rect 1800 -10 1850 5
<< nsubdiff >>
rect -100 1250 -50 1265
rect -100 980 -85 1250
rect -65 980 -50 1250
rect -100 965 -50 980
rect 1800 1250 1850 1265
rect 1800 980 1815 1250
rect 1835 980 1850 1250
rect 1800 965 1850 980
<< psubdiffcont >>
rect -85 545 -65 815
rect 1815 545 1835 815
rect -85 260 -65 380
rect 1815 260 1835 380
rect -85 5 -65 125
rect 1815 5 1835 125
<< nsubdiffcont >>
rect -85 980 -65 1250
rect 1815 980 1835 1250
<< poly >>
rect -100 1305 1550 1320
rect 0 1265 50 1280
rect 100 1265 150 1280
rect 200 1265 250 1305
rect 300 1265 350 1305
rect 400 1265 450 1280
rect 500 1265 550 1280
rect 600 1265 650 1305
rect 700 1265 750 1305
rect 800 1265 850 1280
rect 900 1265 950 1280
rect 1000 1265 1050 1305
rect 1100 1265 1150 1305
rect 1200 1265 1250 1280
rect 1300 1265 1350 1280
rect 1400 1265 1450 1305
rect 1500 1265 1550 1305
rect 1600 1265 1650 1280
rect 1700 1265 1750 1280
rect 0 950 50 965
rect -95 940 50 950
rect -95 920 -85 940
rect -65 935 50 940
rect -65 920 -55 935
rect 100 925 150 965
rect 200 950 250 965
rect 300 950 350 965
rect 400 925 450 965
rect 500 925 550 965
rect 600 950 650 965
rect 700 950 750 965
rect 800 925 850 965
rect 900 925 950 965
rect 1000 950 1050 965
rect 1100 950 1150 965
rect 1200 925 1250 965
rect 1300 925 1350 965
rect 1400 950 1450 965
rect 1500 950 1550 965
rect 1600 925 1650 965
rect 1700 950 1750 965
rect 1700 940 1795 950
rect 1700 935 1765 940
rect -95 910 -55 920
rect 75 910 1650 925
rect 1755 920 1765 935
rect 1785 920 1795 940
rect 1755 910 1795 920
rect 75 905 90 910
rect 30 890 90 905
rect 30 885 45 890
rect -100 870 45 885
rect 120 870 1650 885
rect 0 830 50 845
rect 100 830 150 870
rect 200 830 250 845
rect 300 830 350 845
rect 400 830 450 870
rect 500 830 550 870
rect 600 830 650 845
rect 700 830 750 845
rect 800 830 850 870
rect 900 830 950 870
rect 1000 830 1050 845
rect 1100 830 1150 845
rect 1200 830 1250 870
rect 1300 830 1350 870
rect 1400 830 1450 845
rect 1500 830 1550 845
rect 1600 830 1650 870
rect 1755 875 1795 885
rect 1755 860 1765 875
rect 1700 855 1765 860
rect 1785 855 1795 875
rect 1700 845 1795 855
rect 1700 830 1750 845
rect 0 515 50 530
rect -95 505 50 515
rect -95 485 -85 505
rect -65 500 50 505
rect -65 485 -55 500
rect 100 490 150 530
rect -95 475 -55 485
rect 75 475 150 490
rect 200 505 250 530
rect 200 485 215 505
rect 235 485 250 505
rect 200 475 250 485
rect 300 505 350 530
rect 400 515 450 530
rect 500 515 550 530
rect 300 485 315 505
rect 335 485 350 505
rect 300 475 350 485
rect 600 505 650 530
rect 600 485 615 505
rect 635 485 650 505
rect 600 475 650 485
rect 700 505 750 530
rect 800 515 850 530
rect 900 515 950 530
rect 700 485 715 505
rect 735 485 750 505
rect 700 475 750 485
rect 1000 505 1050 530
rect 1000 485 1015 505
rect 1035 485 1050 505
rect 1000 475 1050 485
rect 1100 505 1150 530
rect 1200 515 1250 530
rect 1300 515 1350 530
rect 1100 485 1115 505
rect 1135 485 1150 505
rect 1100 475 1150 485
rect 1400 505 1450 530
rect 1400 485 1415 505
rect 1435 485 1450 505
rect 1400 475 1450 485
rect 1500 505 1550 530
rect 1600 515 1650 530
rect 1700 515 1750 530
rect 1500 485 1515 505
rect 1535 485 1550 505
rect 1500 475 1550 485
rect 1600 475 1850 490
rect 30 460 90 475
rect 30 450 45 460
rect 1600 450 1650 475
rect -100 435 45 450
rect 120 435 1650 450
rect 0 395 50 410
rect 100 395 150 435
rect 200 395 250 410
rect 300 395 350 410
rect 400 395 450 435
rect 500 395 550 435
rect 600 395 650 410
rect 700 395 750 410
rect 800 395 850 435
rect 900 395 950 435
rect 1000 395 1050 410
rect 1100 395 1150 410
rect 1200 395 1250 435
rect 1300 395 1350 435
rect 1400 395 1450 410
rect 1500 395 1550 410
rect 1600 395 1650 435
rect 1755 440 1795 450
rect 1755 425 1765 440
rect 1700 420 1765 425
rect 1785 420 1795 440
rect 1700 410 1795 420
rect 1700 395 1750 410
rect 0 230 50 245
rect 100 230 150 245
rect -95 220 50 230
rect -95 200 -85 220
rect -65 215 50 220
rect -65 200 -55 215
rect -95 190 -55 200
rect 200 205 250 245
rect 300 205 350 245
rect 400 230 450 245
rect 500 230 550 245
rect 600 205 650 245
rect 700 205 750 245
rect 800 230 850 245
rect 900 230 950 245
rect 1000 205 1050 245
rect 1100 205 1150 245
rect 1200 230 1250 245
rect 1300 230 1350 245
rect 1400 205 1450 245
rect 1500 205 1550 245
rect 1600 230 1650 245
rect 1700 230 1750 245
rect 200 190 1850 205
rect 0 180 50 190
rect 0 160 10 180
rect 30 160 50 180
rect 0 140 50 160
rect 100 140 150 155
rect 200 140 250 155
rect 300 140 350 155
rect 400 140 450 155
rect 500 140 550 155
rect 600 140 650 155
rect 700 140 750 155
rect 800 140 850 155
rect 900 140 950 155
rect 1000 140 1050 155
rect 1100 140 1150 155
rect 1200 140 1250 155
rect 1300 140 1350 155
rect 1400 140 1450 155
rect 1500 140 1550 155
rect 1600 140 1650 155
rect 1700 140 1750 155
rect 0 -25 50 -10
rect 100 -35 150 -10
rect 100 -55 115 -35
rect 135 -55 150 -35
rect 100 -65 150 -55
rect 200 -35 250 -10
rect 200 -55 215 -35
rect 235 -55 250 -35
rect 200 -65 250 -55
rect 300 -35 350 -10
rect 300 -55 315 -35
rect 335 -55 350 -35
rect 300 -65 350 -55
rect 400 -35 450 -10
rect 400 -55 415 -35
rect 435 -55 450 -35
rect 400 -65 450 -55
rect 500 -35 550 -10
rect 500 -55 515 -35
rect 535 -55 550 -35
rect 500 -65 550 -55
rect 600 -35 650 -10
rect 600 -55 615 -35
rect 635 -55 650 -35
rect 600 -65 650 -55
rect 700 -35 750 -10
rect 700 -55 715 -35
rect 735 -55 750 -35
rect 700 -65 750 -55
rect 800 -35 850 -10
rect 800 -55 815 -35
rect 835 -55 850 -35
rect 800 -65 850 -55
rect 900 -35 950 -10
rect 900 -55 915 -35
rect 935 -55 950 -35
rect 900 -65 950 -55
rect 1000 -35 1050 -10
rect 1000 -55 1015 -35
rect 1035 -55 1050 -35
rect 1000 -65 1050 -55
rect 1100 -35 1150 -10
rect 1100 -55 1115 -35
rect 1135 -55 1150 -35
rect 1100 -65 1150 -55
rect 1200 -35 1250 -10
rect 1200 -55 1215 -35
rect 1235 -55 1250 -35
rect 1200 -65 1250 -55
rect 1300 -35 1350 -10
rect 1300 -55 1315 -35
rect 1335 -55 1350 -35
rect 1300 -65 1350 -55
rect 1400 -35 1450 -10
rect 1400 -55 1415 -35
rect 1435 -55 1450 -35
rect 1400 -65 1450 -55
rect 1500 -35 1550 -10
rect 1500 -55 1515 -35
rect 1535 -55 1550 -35
rect 1500 -65 1550 -55
rect 1600 -35 1650 -10
rect 1600 -55 1615 -35
rect 1635 -55 1650 -35
rect 1700 -25 1750 -10
rect 1700 -35 1795 -25
rect 1700 -40 1765 -35
rect 1600 -65 1650 -55
rect 1755 -55 1765 -40
rect 1785 -55 1795 -35
rect 1755 -65 1795 -55
<< polycont >>
rect -85 920 -65 940
rect 1765 920 1785 940
rect 1765 855 1785 875
rect -85 485 -65 505
rect 215 485 235 505
rect 315 485 335 505
rect 615 485 635 505
rect 715 485 735 505
rect 1015 485 1035 505
rect 1115 485 1135 505
rect 1415 485 1435 505
rect 1515 485 1535 505
rect 1765 420 1785 440
rect -85 200 -65 220
rect 10 160 30 180
rect 115 -55 135 -35
rect 215 -55 235 -35
rect 315 -55 335 -35
rect 415 -55 435 -35
rect 515 -55 535 -35
rect 615 -55 635 -35
rect 715 -55 735 -35
rect 815 -55 835 -35
rect 915 -55 935 -35
rect 1015 -55 1035 -35
rect 1115 -55 1135 -35
rect 1215 -55 1235 -35
rect 1315 -55 1335 -35
rect 1415 -55 1435 -35
rect 1515 -55 1535 -35
rect 1615 -55 1635 -35
rect 1765 -55 1785 -35
<< locali >>
rect 455 1280 1850 1320
rect -95 1250 -5 1260
rect -95 980 -85 1250
rect -65 980 -35 1250
rect -15 980 -5 1250
rect -95 970 -5 980
rect 55 1250 95 1260
rect 55 980 65 1250
rect 85 980 95 1250
rect -95 940 -55 970
rect -95 920 -85 940
rect -65 920 -55 940
rect -95 910 -55 920
rect -95 815 -5 825
rect -95 545 -85 815
rect -65 545 -35 815
rect -15 545 -5 815
rect -95 535 -5 545
rect 55 815 95 980
rect 55 545 65 815
rect 85 545 95 815
rect -95 505 -55 535
rect -95 485 -85 505
rect -65 485 -55 505
rect -95 475 -55 485
rect 55 515 95 545
rect 155 1250 195 1260
rect 155 980 165 1250
rect 185 980 195 1250
rect 155 585 195 980
rect 255 1250 295 1260
rect 255 980 265 1250
rect 285 980 295 1250
rect 255 970 295 980
rect 355 1250 395 1260
rect 355 980 365 1250
rect 385 980 395 1250
rect 155 545 165 585
rect 185 545 195 585
rect 155 535 195 545
rect 255 815 295 825
rect 255 545 265 815
rect 285 545 295 815
rect 255 535 295 545
rect 355 585 395 980
rect 355 545 365 585
rect 385 545 395 585
rect 355 535 395 545
rect 455 1250 495 1280
rect 455 980 465 1250
rect 485 980 495 1250
rect 455 815 495 980
rect 455 545 465 815
rect 485 545 495 815
rect 455 535 495 545
rect 555 1250 595 1260
rect 555 980 565 1250
rect 585 980 595 1250
rect 555 585 595 980
rect 655 1250 695 1260
rect 655 980 665 1250
rect 685 980 695 1250
rect 655 970 695 980
rect 755 1250 795 1260
rect 755 980 765 1250
rect 785 980 795 1250
rect 555 545 565 585
rect 585 545 595 585
rect 555 535 595 545
rect 655 815 695 825
rect 655 545 665 815
rect 685 545 695 815
rect 655 535 695 545
rect 755 585 795 980
rect 755 545 765 585
rect 785 545 795 585
rect 755 535 795 545
rect 855 1250 895 1260
rect 855 980 865 1250
rect 885 980 895 1250
rect 855 815 895 980
rect 855 545 865 815
rect 885 545 895 815
rect 855 515 895 545
rect 955 1250 995 1260
rect 955 980 965 1250
rect 985 980 995 1250
rect 955 585 995 980
rect 1055 1250 1095 1260
rect 1055 980 1065 1250
rect 1085 980 1095 1250
rect 1055 970 1095 980
rect 1155 1250 1195 1260
rect 1155 980 1165 1250
rect 1185 980 1195 1250
rect 955 545 965 585
rect 985 545 995 585
rect 955 535 995 545
rect 1055 815 1095 825
rect 1055 545 1065 815
rect 1085 545 1095 815
rect 1055 535 1095 545
rect 1155 585 1195 980
rect 1155 545 1165 585
rect 1185 545 1195 585
rect 1155 535 1195 545
rect 1255 1250 1295 1280
rect 1255 980 1265 1250
rect 1285 980 1295 1250
rect 1255 815 1295 980
rect 1255 545 1265 815
rect 1285 545 1295 815
rect 1255 535 1295 545
rect 1355 1250 1395 1260
rect 1355 980 1365 1250
rect 1385 980 1395 1250
rect 1355 585 1395 980
rect 1455 1250 1495 1260
rect 1455 980 1465 1250
rect 1485 980 1495 1250
rect 1455 970 1495 980
rect 1555 1250 1595 1260
rect 1555 980 1565 1250
rect 1585 980 1595 1250
rect 1355 545 1365 585
rect 1385 545 1395 585
rect 1355 535 1395 545
rect 1455 815 1495 825
rect 1455 545 1465 815
rect 1485 545 1495 815
rect 1455 535 1495 545
rect 1555 585 1595 980
rect 1555 545 1565 585
rect 1585 545 1595 585
rect 1555 535 1595 545
rect 1655 1250 1695 1260
rect 1655 980 1665 1250
rect 1685 980 1695 1250
rect 1655 815 1695 980
rect 1755 1250 1845 1260
rect 1755 980 1765 1250
rect 1785 980 1815 1250
rect 1835 980 1845 1250
rect 1755 970 1845 980
rect 1755 940 1795 970
rect 1755 920 1765 940
rect 1785 920 1795 940
rect 1755 910 1795 920
rect 1655 545 1665 815
rect 1685 545 1695 815
rect 1655 515 1695 545
rect 1755 875 1795 885
rect 1755 855 1765 875
rect 1785 855 1795 875
rect 1755 825 1795 855
rect 1755 815 1845 825
rect 1755 545 1765 815
rect 1785 545 1815 815
rect 1835 545 1845 815
rect 1755 535 1845 545
rect 55 505 1695 515
rect 55 485 215 505
rect 235 485 315 505
rect 335 485 615 505
rect 635 485 715 505
rect 735 485 1015 505
rect 1035 485 1115 505
rect 1135 485 1415 505
rect 1435 485 1515 505
rect 1535 485 1695 505
rect 55 475 1695 485
rect 55 440 1695 450
rect 55 420 155 440
rect 195 420 755 440
rect 795 420 955 440
rect 995 420 1555 440
rect 1595 420 1695 440
rect 55 410 1695 420
rect -95 380 -5 390
rect -95 260 -85 380
rect -65 260 -35 380
rect -15 260 -5 380
rect -95 250 -5 260
rect 55 380 95 410
rect 55 260 65 380
rect 85 260 95 380
rect 55 250 95 260
rect 155 380 195 390
rect 155 260 165 380
rect 185 260 195 380
rect -95 220 -55 250
rect -95 200 -85 220
rect -65 200 -55 220
rect -95 190 -55 200
rect 155 220 195 260
rect 255 380 295 390
rect 255 260 265 380
rect 285 260 295 380
rect 255 250 295 260
rect 355 380 395 390
rect 355 260 365 380
rect 385 260 395 380
rect 355 220 395 260
rect 455 380 495 410
rect 455 260 465 380
rect 485 260 495 380
rect 455 250 495 260
rect 555 380 595 390
rect 555 260 565 380
rect 585 260 595 380
rect 555 220 595 260
rect 655 380 695 390
rect 655 260 665 380
rect 685 260 695 380
rect 655 250 695 260
rect 755 380 795 390
rect 755 260 765 380
rect 785 260 795 380
rect 755 220 795 260
rect 855 380 895 410
rect 855 260 865 380
rect 885 260 895 380
rect 855 250 895 260
rect 955 380 995 390
rect 955 260 965 380
rect 985 260 995 380
rect 955 220 995 260
rect 1055 380 1095 390
rect 1055 260 1065 380
rect 1085 260 1095 380
rect 1055 250 1095 260
rect 1155 380 1195 390
rect 1155 260 1165 380
rect 1185 260 1195 380
rect 1155 220 1195 260
rect 1255 380 1295 410
rect 1255 260 1265 380
rect 1285 260 1295 380
rect 1255 250 1295 260
rect 1355 380 1395 390
rect 1355 260 1365 380
rect 1385 260 1395 380
rect 1355 220 1395 260
rect 1455 380 1495 390
rect 1455 260 1465 380
rect 1485 260 1495 380
rect 1455 250 1495 260
rect 1555 380 1595 390
rect 1555 260 1565 380
rect 1585 260 1595 380
rect 1555 220 1595 260
rect 1655 380 1695 410
rect 1655 260 1665 380
rect 1685 260 1695 380
rect 1655 250 1695 260
rect 1755 440 1795 450
rect 1755 420 1765 440
rect 1785 420 1795 440
rect 1755 390 1795 420
rect 1755 380 1845 390
rect 1755 260 1765 380
rect 1785 260 1815 380
rect 1835 260 1845 380
rect 1755 250 1845 260
rect -35 180 40 190
rect 155 180 1595 220
rect -35 160 10 180
rect 30 160 40 180
rect -35 150 40 160
rect -35 135 -5 150
rect -95 125 -5 135
rect -95 5 -85 125
rect -65 5 -35 125
rect -15 5 -5 125
rect -95 -5 -5 5
rect 55 125 95 135
rect 55 5 65 125
rect 85 5 95 125
rect 55 -25 95 5
rect 155 125 195 135
rect 155 5 165 125
rect 185 5 195 125
rect 155 -5 195 5
rect 255 125 295 180
rect 255 5 265 125
rect 285 5 295 125
rect 255 -5 295 5
rect 355 125 395 135
rect 355 5 365 125
rect 385 5 395 125
rect 355 -5 395 5
rect 455 125 495 135
rect 455 5 465 125
rect 485 5 495 125
rect 455 -25 495 5
rect 555 125 595 135
rect 555 5 565 125
rect 585 5 595 125
rect 555 -5 595 5
rect 655 125 695 180
rect 655 5 665 125
rect 685 5 695 125
rect 655 -5 695 5
rect 755 125 795 135
rect 755 5 765 125
rect 785 5 795 125
rect 755 -5 795 5
rect 855 125 895 135
rect 855 5 865 125
rect 885 5 895 125
rect 855 -25 895 5
rect 955 125 995 135
rect 955 5 965 125
rect 985 5 995 125
rect 955 -5 995 5
rect 1055 125 1095 180
rect 1455 175 1595 180
rect 1055 5 1065 125
rect 1085 5 1095 125
rect 1055 -5 1095 5
rect 1155 125 1195 135
rect 1155 5 1165 125
rect 1185 5 1195 125
rect 1155 -5 1195 5
rect 1255 125 1295 135
rect 1255 5 1265 125
rect 1285 5 1295 125
rect 1255 -25 1295 5
rect 1355 125 1395 135
rect 1355 5 1365 125
rect 1385 5 1395 125
rect 1355 -5 1395 5
rect 1455 125 1495 175
rect 1455 5 1465 125
rect 1485 5 1495 125
rect 1455 -5 1495 5
rect 1555 125 1595 135
rect 1555 5 1565 125
rect 1585 5 1595 125
rect 1555 -5 1595 5
rect 1655 125 1695 135
rect 1655 5 1665 125
rect 1685 5 1695 125
rect 1655 -25 1695 5
rect -100 -35 1695 -25
rect -100 -55 115 -35
rect 135 -55 215 -35
rect 235 -55 315 -35
rect 335 -55 415 -35
rect 435 -55 515 -35
rect 535 -55 615 -35
rect 635 -55 715 -35
rect 735 -55 815 -35
rect 835 -55 915 -35
rect 935 -55 1015 -35
rect 1035 -55 1115 -35
rect 1135 -55 1215 -35
rect 1235 -55 1315 -35
rect 1335 -55 1415 -35
rect 1435 -55 1515 -35
rect 1535 -55 1615 -35
rect 1635 -55 1695 -35
rect -100 -65 1695 -55
rect 1755 125 1845 135
rect 1755 5 1765 125
rect 1785 5 1815 125
rect 1835 5 1845 125
rect 1755 -5 1845 5
rect 1755 -35 1795 -5
rect 1755 -55 1765 -35
rect 1785 -55 1795 -35
rect 1755 -65 1795 -55
<< viali >>
rect -85 980 -65 1250
rect -35 980 -15 1250
rect -85 545 -65 815
rect -35 545 -15 815
rect 265 980 285 1250
rect 165 545 185 585
rect 265 545 285 815
rect 365 545 385 585
rect 665 980 685 1250
rect 565 545 585 585
rect 665 545 685 815
rect 765 545 785 585
rect 1065 980 1085 1250
rect 965 545 985 585
rect 1065 545 1085 815
rect 1165 545 1185 585
rect 1465 980 1485 1250
rect 1365 545 1385 585
rect 1465 545 1485 815
rect 1565 545 1585 585
rect 1765 980 1785 1250
rect 1815 980 1835 1250
rect 1765 545 1785 815
rect 1815 545 1835 815
rect 155 420 195 440
rect 755 420 795 440
rect 955 420 995 440
rect 1555 420 1595 440
rect -85 260 -65 380
rect -35 260 -15 380
rect 265 260 285 380
rect 665 260 685 380
rect 1065 260 1085 380
rect 1465 260 1485 380
rect 1765 260 1785 380
rect 1815 260 1835 380
rect -85 5 -65 125
rect -35 5 -15 125
rect 165 5 185 125
rect 365 5 385 125
rect 565 5 585 125
rect 765 5 785 125
rect 965 5 985 125
rect 1165 5 1185 125
rect 1365 5 1385 125
rect 1565 5 1585 125
rect 1765 5 1785 125
rect 1815 5 1835 125
<< metal1 >>
rect -100 1250 1850 1260
rect -100 980 -85 1250
rect -65 980 -35 1250
rect -15 980 265 1250
rect 285 980 665 1250
rect 685 980 1065 1250
rect 1085 980 1465 1250
rect 1485 980 1765 1250
rect 1785 980 1815 1250
rect 1835 980 1850 1250
rect -100 970 1850 980
rect -100 815 1850 825
rect -100 545 -85 815
rect -65 545 -35 815
rect -15 615 265 815
rect -15 545 120 615
rect -100 535 120 545
rect 155 585 195 595
rect 155 545 165 585
rect 185 545 195 585
rect -100 380 -5 535
rect 155 450 195 545
rect 220 545 265 615
rect 285 615 665 815
rect 285 545 325 615
rect 220 535 325 545
rect 355 585 395 595
rect 355 545 365 585
rect 385 545 395 585
rect 145 440 205 450
rect 145 420 155 440
rect 195 420 205 440
rect 145 410 205 420
rect 355 390 395 545
rect 555 585 595 595
rect 555 545 565 585
rect 585 545 595 585
rect 555 390 595 545
rect 625 545 665 615
rect 685 615 1065 815
rect 685 545 725 615
rect 625 535 725 545
rect 755 585 795 595
rect 755 545 765 585
rect 785 545 795 585
rect 755 450 795 545
rect 955 585 995 595
rect 955 545 965 585
rect 985 545 995 585
rect 955 450 995 545
rect 1025 545 1065 615
rect 1085 615 1465 815
rect 1085 545 1125 615
rect 1025 535 1125 545
rect 1155 585 1195 595
rect 1155 545 1165 585
rect 1185 545 1195 585
rect 745 440 805 450
rect 745 420 755 440
rect 795 420 805 440
rect 745 410 805 420
rect 945 440 1005 450
rect 945 420 955 440
rect 995 420 1005 440
rect 945 410 1005 420
rect 1155 390 1195 545
rect 1355 585 1395 595
rect 1355 545 1365 585
rect 1385 545 1395 585
rect 1355 390 1395 545
rect 1425 545 1465 615
rect 1485 615 1765 815
rect 1485 545 1525 615
rect 1425 535 1525 545
rect 1555 585 1595 595
rect 1555 545 1565 585
rect 1585 545 1595 585
rect 1555 450 1595 545
rect 1625 545 1765 615
rect 1785 545 1815 815
rect 1835 545 1850 815
rect 1625 535 1850 545
rect 1545 440 1605 450
rect 1545 420 1555 440
rect 1595 420 1605 440
rect 1545 410 1605 420
rect -100 260 -85 380
rect -65 260 -35 380
rect -15 260 -5 380
rect -100 135 -5 260
rect 255 380 1495 390
rect 255 260 265 380
rect 285 260 665 380
rect 685 260 1065 380
rect 1085 260 1465 380
rect 1485 260 1495 380
rect 255 250 1495 260
rect 1755 380 1850 535
rect 1755 260 1765 380
rect 1785 260 1815 380
rect 1835 260 1850 380
rect 1755 135 1850 260
rect -100 125 1850 135
rect -100 5 -85 125
rect -65 5 -35 125
rect -15 5 165 125
rect 185 5 365 125
rect 385 5 565 125
rect 585 5 765 125
rect 785 5 965 125
rect 985 5 1165 125
rect 1185 5 1365 125
rect 1385 5 1565 125
rect 1585 5 1765 125
rect 1785 5 1815 125
rect 1835 5 1850 125
rect -100 -5 1850 5
<< labels >>
rlabel metal1 -100 680 -100 680 7 VN
port 3 w
rlabel metal1 -100 1115 -100 1115 7 VP
port 5 w
rlabel locali 1850 1300 1850 1300 3 Vout
port 7 e
rlabel poly -100 1310 -100 1310 7 Vbp
port 6 w
rlabel locali -100 -45 -100 -45 7 Vbn
port 1 w
rlabel poly -100 445 -100 445 7 Vcn
port 2 w
rlabel poly -100 875 -100 875 7 Vcp
port 4 w
rlabel poly 1850 485 1850 485 3 V1
port 8 e
rlabel poly 1850 195 1850 195 3 V2
port 9 e
<< end >>
